PK   Ci�St��R$  k    cirkitFile.json��n$Ǒ�_E��b2�P���%X�a/,�7�P��L,E�6IɆ�ڗ�gڌ����՝5��J�f.D���ʎ�Ȫ���j��0�5��nl~w7�wWo�]_���?�/��^_���k��v�\����n��n4�nl��>�i��#��7�RkB��T��L1�.Nվ���z�ͷ��@bې�A�`'f�*�Ƌ�
�	b��m��A�`�B� U�M)f�*ئ3��������ƻǦrU�Қ��Ʉ0���Z2E�zJҝK_K{%���R���AV,�( a�$גj�$y�K$
/��2hz�'�OPI?���Aڋ�������N寧����~z�]�J�'��O �����J�����"�mU,1ăv�}���b����)���.�-̡MҥI��v����'Ob�9)����'Pb��n-���{'��b�y�)���lo_}�?B@6�=��C�C�X"Q�C���|�`ԋB~���D�y�;���1��B~�𢬆��Q/�ۈ%��n#�H�X"Q��6b�"��X"Q�ob�D!�]�%��!�X"Q s��n��]�D���N�D���N�D���N�D���N��m�<v�%�<v�%�<v�%�<v�%�<v�%�!�<vFy�K$
y�K$
y�K$
y�Kئ��N�D���N�D���΅Ļ�ǝٵ7���yw��n��? ����r��#,]Jϱ��;(a�l��9�wP:����c��X�t��K9ֻ��JGX�4��z��A�K���X�
�wP:��٦�zWb�����6ֻ
����t�����X�t���w{��cpf��#0����]��p~A������|��?p���#0�K��i`���o���gX>����`�����|�6=�?pց�#0����y`���+	����,��xx��`��������,��x�	�?��#p������X>������G`>^-��`��������,��x��?p���#0�-��?�|��Uq�|�6�by��\����`�x��p��#0�B�N]�|����`������|�z��-�Z��ŃSN]�|��e�`������|�h�8u���������.X>��Be����G`>^b��`��ǋñ�p���#0/k��?�|���`������|\J �8������ ��C/A���p���#0� ��?�|��`������|\��8�����˔���X>�q���`��ǥa����,�����?p���#0����?�|��BB`������|\	�z�:z�:8����#��,�����?p���#0���?�|��R_`������|\��_�?�|���j`������|\�8������/�W�Zq]�������EH7��n!��5ߗg��M�_�������������:76?����K�¯ 9Q/��L���KO�D�?�໵�q�ݭ�]����ݮd�;�����D��;�&>�'���$��N���O�O/��(�8��w��Sr�(��T�N_HO_�N_JO/����g��^��Um�
��^�/irC�ǲO�ce�PG��Cm����܈?����˖z�b�Fn�Sw�5d��,�~�E<s����g��}oc�b0��*ӵeeZ��/����3g�j�~�1����Xv�	}��ܐ>�`�����Μ=������Yo�0�&L]a�2:3���T��t>��z���|=U�j�>L�j�>J�j�>��j����]��~��^�q��~��������bl����	>����[U.����4����4?��i�n^V�u��bL�:�J�M(��t~�L�Ot]����>{V��Ϟ�|��g5?3�S���L]�hB]���n�q�\��G:{��h��٭O��ZccL�7DS�љ�������Ey��Y���<�o����~w��'ɰ%]���$;^Jh�=����	IHh������iSHh�J����UHh������y_�,�����GQ�"	�g�A!�qa��T}U!d�n��~j��w_}��h��	��s�W�2�J5}i����i��u��.d:����?D!S��v�/E1�J�kw���h�rz�`��R�y�
i,��q���Ih`	���QJ��" �����}��OJ�~������2�⸃�QJ�g* &�8���(���,�;XG)�Ӏ�`q�������Ka:���QJ\��4+���Ǚ�î,�{XG)q�*S�;^�Ͻ�	�QJ\g	����QJ\���6G)q�,�XG)q}nN7)���QJ\[����QJ\����QJ\� ���#,���xM=�	�#,���x�7�	�t�x�#,���x�/�	�#,���x}*�	�XG)�:J,��8���}!���Z����J*���j��e�pU�����j���pU�����j��2ApU�����._��a�`%�4R�����VRaMc_��a�`%V��!��}�`%V��'��}�`%V��-��}�`%V~'X'1�ɸThI���m��V)�RJ�t�.�I�H'�R�%Z~�\�[��K��th��you20Zҡ�w�u����ThI���0�x����В-����V'S�%Z^S��NF�BK:��6F�[��L��thy��΃��L��thy����:y�
-���+o���)=��˜N^�t�2Zҡ�5p:���e*��C�k�t����ThI���$�x����В-����V'/S�%Z^#��N^�BK:��b�o煊PY��:y�
-���y1I'/S�%Z^{��N^�BK:���Z�[��L��thy-���Jo+*�����y�����e*��C�k�u����ThI��k�x����В-�J��V'/S�%Z����N^�BK:�\�B�[��L��th����A'/S�%Z�%��N^�BK:�\E�[��L��th�����:y�
-��r�o�V�)-%��˂N^t�2Zҡ�A:���e*��C˵�t����ThI��k8�x����В-ע��V'/S�%Z����m���ThI��k��x����В-�8��V'/S�%Z�զ�N^�BK:�\sN�[��L��th�v���JU>��|��eQ'/�:y�
-��r-Cou�2Zҡ嚌:���e*��C˵%u����ThI��kd�x[��e*��C˵>u����ThI��k��x�����R��]���f*h2!�i��LQ����;����F��ڴUV��nTY��Qe�����g��a�!�Ju�*+��7��T�ި�R�yk�u^L��o��ܨh����{Um�Y)�Uf���VL^�st�̡o�U�Ћ�w���^��zz��܋�;Ln��o���Bu��!
Ufe��2�^|���V��}��̽x�W�V�C/>ކy�L��P�;Lo��bb���/dJ�ܐG�X�I&V�
u4޻>�v�k3F59*Yʖz�b�H��*]0u�[C��ˢ�G_��,Y*Yu}���ءL��tmY�և~��a���2K��E�1����Xv�	}�.��>�`�����.�d�\dl�
g�)�T�0u������C�]7tS�'�R�8~�R�8~�R�x��R�x��R�x��R�8f̻��]���a�a���1�X��ض�),9|����[U.�ө�4f|�sT.����f�\��/�t7	���{��3��*�nk]�ap}�/Y*}�R��K���T�tQ?���ф�"S�3E�&W�!��rn�*}�>�?Bh���5���at��i�z7�}Q^f�Ry���,�<�7���x�������a����q�޾�۾uHh?�!	� D ����$��ނ���Se"��~�B�O�A�@B��@Hh?�!	�)1!�qa�	�QJ��X,v,x����&X�&X G)f�1L�N� �R:̭c�`q���8J�0�a�qpXw�8�R:<��0�⸃�q����	�,����0L�8�`q�txT�I�aq���8J�����p3)��X��8�R�b\0&X��8�R��O0&X��8�R�bC0&X�8�R��60&X�8�R�b*0&ܜ8nR�,������	�,������	�,���xQ?��,�GXG)�"r,�GXG)�e��&��&,�GXG)��R,�GXG)�bF,��8�R��s0&X/`q|Mi�B��BK��~�@�TXI��6�E�hU�����j��K�*�WVRa�͢�Z�+����K��E�����A*�.j�@�`%�4FQ�uQ��+���fQ��
�U��TXm�(p�V���J*��Y�A�}�`%V~'X'1�ɸThI���m��V)�RJ�t�.�I�H'�R�%Z~�\�[��K��th��you20Zҡ�w�u����ThI���0�x����В-����V'S�%Z^S��NF�BK:��6F�[��L��thy��΃��L��thy����:y�
-���+o���)=��˜N^�t�2Zҡ�5p:���e*��C�k�t����ThI���$�x����В-����V'/S�%Z^#��N^�BK:���U�[��L��thyͮ΋I:y�
-����cou�2Zҡ�5�:���e*��C�k�u�Uz[Q�uE�����e^'/S�%Z^���N^�BK:�\c@�[��L��th�V���:y�
-��r�ou�2Zҡ��:���e*��C�58T�:y�
-��r-ou�2Zҡ�(:���e*��C˵]t����ThI��k��x���Li)�N^t򲠓��В-���V'/S�%Z�}��N^�BK:�\�I�[��L��th����:y�
-��rM-o�N^�BK:�\L�[��L��th�ƙ��:y�
-��r�6ou�2Zҡ�s:���e*��C˵�t�U��T�C'/�:yY���ThI��k�x����В-�d��V'/S�%Z�-��N^�BK:�\#S��B'/S�%Z����N^�BK:�\�T�[��L���h_l[�0��5SA�	ahM;�d��U���ع��7��Ԧݨ�RMv��J�*+��7����ި�R�z��J=�*+�7���|���@��{�6}�*��k[�n����L��`���6�[e0�xm3έ2����k�Tn���⵽ ��`z�ڎ�[e0�xm_íw]L/^�=��LI����>���T���{ׇڎ�smƨ&G�"K�R�\LiY���zk�uYt��x�%K�"K���{;;�	]W��-+���}9Lu5\f�R��2�6x��n4��ҥ��lp��uߖ�e�,��,��U�7E�j��0u�}H=��n��DY*Cg���ș�r1pf�\��Y*�]���8�w�/v�<P��t��c�<���f��bl����	>�Tc썭*����G3��9*��L��E�T.��c����P�	Eՙ�O�I����0�>×,���d�\�%K�� �tQ?���ф�"S�3E�&W�!��rn�*}�>�?Bh���5���at��i�z7�}Q^f�Ry���u��&C�o�w���ϫ�T]_�x��w�m?��]s�����o��p��;��/�h ����Q6�����ʥ������k/7_t��拮}!>})�NE�'��Ӌ������wO�DSQ®�Da���lMxzѥ��Ͼyn_������xI7F��D{+�^�-� /	�)����!�n����4&l�S��oh��O??�����Ϗ����
i����f��tO����-�P�;5�BܩQ�q�TƯ ����҉�_A�)P�i���;`6C!��PH�F �)H�ϔ`��t�B!�7�U<>������L�AB�t�M��&� AD<熡O�%��t§�����}�޾���4������f�z���{~��H.�%���)�����b��r!�Xb��@H!��/WR�%���b��r	!�Xb��BH��՟�C��P�J,qX�!�b�`�����HV��r��z{�G���GT�����Bʸ�tB�����XJ�ƨ���^�r��X��N��NˠnK! ��5ˡ��B@Xw��.�8,Ȓr�ew��X'�z-��uH�5+Τ������5oR@�u��+�8���r ��l�h$�u{@����+��}� ��K�a�<�j����W��;8��d�= �5x�  {@,�k�F* @,���\�7� p �o _�o� �@�#&��5 «\���8 �4 �\���8 �4 �\���g �i�S��p �i�S�7p ��!��i�S��p �i�S�.p �i��r.�	� ��O��_uZI���L���G`>�,
��� �a��g�E�S��?,��l��h���G`��o��[�"!��X>��ؿ�N�ϋ�#0_��[�!��X>��f��N����|�Yl�Ӄ���#0�m8�� �a���/b���LHhB~��!<��!�<�Љ�30!�	�m]���lLHhB~��!:#��_|F{��J���&�ײ��30!�	�r����LHhB~��!:C����G{��R���&��jt�&$4!��@{��S���&�h�OL��L�y�C�)���		M�ke���0!�	y��Ct�&$4!�QB{��S���&��Uh�y
��Є�6�!:O�pYvi�����1���0!/�C��N[���&���h�i��Є��!:m��n�=������xt���i��Є�B�!:m����=D�-`BB�Rd���LHhB^F�����		M�K����0!�	y�:�À�S���&��h�y
��Є\6 �!:O��K�=D�)`BBr�����)�)�<%���S���&�2h�y
��Є\��!:O��˓�=D�)`BBri���<LHhB.�0��0!�	���Ct�&$4!��A{��S���&�RBh�y
��Є\	�!:O��K8�=�/����G�)��Dt�&$4!��B{��S���&�_h�y
��Є\��!:O��˭�=,�y
��Є\*�!:O���ܡ=D�)`B�D�q��E�í{T
�/Jnl�(��y���l���K��K7�_��~Q tc�Eaϭ�K�=���Nl�!���/�$[�Ӣ��V�Eqޭ�N�ܷl�&��w�ھ�����I~~���۽���j�މ�J�޲����o�ޥ����eP�t��ܪwbo@�]ĝ�~�����a%ߏ�L[�E��&7�aT?�}���B�����ڳ����g�_��;�Fn�Sw�5d��,�~�E<w���g�������`B�U�k�ʴ>�C_S]�Ο�������b0cٍ&�]��C���w���r:w���g�?�X�zS��6a�
S�љчԷ�n観�Y�όb�ڟ�f�?3�jf����<���qb��;Ӂ��=H���o8�	ƪ,ƶM��|���[U.E���4���?rڟq0���bL1<�J�M(��t~�L��t]���g?V�3�?���ϟ��\*\���L]�hB]��ߙ"N����H�o���|~��]<���[�MFg*�ƮwS���g�ߟ����n���I�Wo��K\����2<>�1��xl��M��so�I�<����y�`N����׉��q�-ܬ�-�p��q�-�p��q�-����tڌ���� g��Aν�U����9�����<o;�d���Ns�_'�|1^�ӓ_4H��i߉��G��M:�2ǣ������#���+�Ւ��D���:A�D���<A�D���8A�D�i�x�(��H؏�	�BJ$�G�Q)%�L��ْ�9�t�����D��D$��\�Z6Ź$��ljD�Ȟ z�7?�=<������o/�R�M�O�-���f�#K"i���G5����q��cs�v�-Î��.?�Q��:��!w8䖇��_
�Cay(���p�X*����p�Z����!zv��v�{;�~г�4����#��--�gK���k���6/z���t���<<r7��R�o\���ؘҽ�_�	������ln�鑻�/q��������ß������q�x3�)�����=�Q����w���w>z}�C{���|�G܁��n�U��������/���۩�}���q������v|�o��nvcJ���H����ij�ǧݸ;���^�솧��{ IBI�����>����ѿ)�?������&�{j�r���!e�eL�uloZ�.Y���/e,C��{s������6Y�W���t��=��ӻ�O�ͮ�0���:1l�&������{��+�u*���z���V�kM�����J�WZP�֢Xi\�<-��!:��p��/~�W��/E��$����b�[kaWZ�z���"<�G>��G������<X\�Á��y>��<���|;�����ǧ������a��7���~*��u|���^D������������g�����sS8\���������;���u��R]�R`�k�����o��1M������>���{
�8<�sBo��O������������".�🟾���g�>�C{7<��;���� �u�.��z�
��m�u����[�>E�X��m��a,M�m4#�)�����."oΜiN䝿{���7/�5�G>���Lo����^��>�I�n��}��������+�S���g�fz�����Oqb w�MY]�G�'#�S�>���No�G�9��K{s�S���|0�?���P}4>���M�U�a(Fq6�����gE��tg��P�.}��ޤ�6���H�-��=�z�50��:��Ii
^�G���6G��x��5����#Ν�U|Փ܇�>�H'��CK�ӿw�N����
}[&���o_!~��4lq��髯�E_��|����0��Q���~�>}[,_���?���TUL_
?���tu�3�R��v*�8N]]����bCη�����8�4s_��Y���
Ͽ��#�;�oJW�1�Xt�Jڑ�^t��H~����{}[J�߸���.���'~m��i ����Q�(�u����?nb(�ŭ�/��h�TL}}���E�OF��GIc�O���ҙ���{��"��3ө��Ǿ���?�PK   Ci�S%�$�& �\ /   images/66379bcf-d80b-4bdc-b204-78d4e16074e1.png�|�?����A�0RʦT���2
�H6%�}�M��lIFd��"d��2#�K9F��ut�c�^ϣ�z���>�n��<��c\�u���	��V��Ƕ�B�]��r��_�BQ}�CW~\����]n�/���{n���{].��P\���w���"����������Wk�����'{7�.�Bή��y6�(��9}�糃&���HK�B
$����X����$�Ҧ-�7t�T2L�ZU�sn��xx�뮋�Z���;xKq��F����(>�{ʔ��]޿�}�6t��L��C���:��#k��v�+�$:�����-3� �x1�y���?�ϭ�y�y�����v[�)zs�~�?#�~���n���n�*�7��F	���3`#( � //�o�n�m�%X���k�c�j�k�K77H5���z%���L����#�`S�3jW��'��:#��چ��̛��MR��&��9��!�׿N�=V�k^��;p���\�$��+�]�����\[/\���^ޞJPxX��π�
��G{a������Z�~��Z�
���H����q�����q�v��p@�����alj� ����Z��nT�����&��@Eŕ��۳�f�z-㿗�S�`����J[�^�܆�nL|,�Z�����i\zp�k����CAۛi��i^i˽�����p���F��x�b�|�ֻZ��8i���f��z��9W�Y��������a\�[��6>�m�"sl<��#�{|���*h�2�4���=��^��5�lv�lF׮�׮E�mk�g��Éh��W�>(�����ʰ�_0���^0g_��MT
���O��و=�\�}������9J��]��]���}�?�4>����y���g�{�o��[����.z������

	5���ܼs������7��E�}noWM���6�et$����������c&}�;)@%��i:u||�������8l;��v��4�p���|�EZj�
�cɷs�3�wF5���
�?��a�w�z�.Ǆ��3MbӢ����8I�yz���<��*��I��}��у��0��3
��ϑ�݁�*�W]M+=�y���|.�%ԑ"�\X�l���մ��9;;�7K�R~��S2�G\���OH���-~��G~�GJ�����������OL�CL1��p!b��\�щ����}N�U1119�~r����Mm�Bukdt�TWW�,�/�B�̚���o�.�5�r��VAAJK,��ZX*����2���=��_b�o��(��fs�?c�l�~@`�V����W 7kqۼ��?-����kr��R��;?B/�cyn =������j��U�Qv�NNBC�Ai/���������7����RC���}���h�DF+�]�ئodh�,�=���ޢ�[4�݆��#�k��������9��*�sm3W配�d	�tS�z|�&4̡t� Iޓ)^7�:�O��ma��w�}oA��򗝷3�v�R�Q���ѥ��H	���5�n��L�$�����2*�&��6��6���@_���d��I���"4|�ru�J"�`�Q�`�C*]u�e�m�[��b��*���\��[`��@��&��,��P�s���@&����E����u+���S��#٥F�z-tv�`e?�yZ�n���gv[��#�*�3�x���F�X�j�|��kc��櫥�&S߭C(R�ZRк�h�SUU�gjp�t�9z�mc�i�˝Gc�b|~&F�G�A/��+0%�j�@��zG�#�������w����jf�P=��ÙV�*a	'`�R�r�~�}?���.��~��M��( $�͕u�z����-������9�𥱎K+�{��p�.��cBa���������ֻ��M�7�T�tWX �o�ø�+k�1����ٖ��&�~�
��4�T��GBQi���	��h%����Lr�iM���߯Т� ����*��4���	�(a����nj�1���Ĺ��RZc��I6f�䯩.4�0(�1��?Z�~�=[�V>(��ԗ)8�Ǖ&}���z���l(�"�<��(6ÊW�)E��U	��|��i �@�,�(3#��p[�;�R��n
a~��2�e�`�^�S�HԀ�
����Ai\i���^V�W��Ǉp#Dje��P$QC�:��&��e��΀�I�K0޽��3�����H�K!�a8
�J�Z�q�mvRK�lbZZ4�D
��BYy��0��J[G�[�����L� �(��� �JD{qq�"��S.U!dz�/�k(�9Vo�ͤ�~jx��?���hjj�x�~*WLt�;kʍ���z $*��(T?�?wha��)���Z�ת���~l&�W�����OÄ�R���PQ9f�>��	��9�\����Y�"�Exޒ����g����33-�9x�FA&���Oa�\��*ZؔB��ۨ�y8
�Ee���{2%<�%K�lP�"0��a�eI	KL��Z�Ps��n擰}��k�����$�XM~}c"����K����|/X~���@�b���Ѐ��x�R{M���y��Mv���)���/�|#B�UT��f\T�������c��E����<�6|�o���T�U�J@���K����^+�����`>Cs�#�0 ��#�* ��d�X~ZA�pn�|8f�̂����Q����I��װ#g0�������a84.���Q�j%q6�#�/{��)A�B[�I��ڴn�:[�1�+�P�%@�����tƢ�8y�VpZC�W�x�����4��!5q�"d�&�?x�;Cd7B�PC���|J	�s� ��܋eB�1z�?`ƫ�c*S� �c20��BWiEx��U����<��!�+����0��0ً�4%n2�Q{w�A�"��B��kf��/�QøT�84��˕Z����v���M�.�=qm�t_eA�MNN��1?_;��� ��65��/�_�Mў�����L"etM!Ka���P�k�</�F'��4�iK�yYǥL�?�Y�~�&��2>���ixڊ?)����v�	q�ȗ�P���O�ׯ��`�M	+84R�nS2E�f���~fv�����LԨD�\��1<�s
P�ׅQ3�-*b�6��]6��ٙ|yD]�/�[��4��GG�FxmZ4�������p�TW�^���(��J3��D4�W�vv��AJ�P;L��C)���+"#�>��Hloo��Y	0"Q�]x��A�F����>��e�h���=�V|[2��W.^�?ă]442"���u3/��~�y���ط�}Gs��%t��8[��`[�6k#d�����߈<�-�>.�ȠH�����'�E��	�>���^TS�
��i�t��t�^X__/*)�E.��-C����w�[����h��K�T��obn����m%R/ �ʭu*�	eW��ѱ���I����F4K���P��%��c0��NR�)>X��xV�� �z�"K���9]��@���e�Z�!�Ջ>O�w�#S��%z]a�4
o.( �7`W(*Q�\�����6]3b|��}pJ��i�o#��S������deeÖ����d ��3K�w!�;%%�|y�s :	%���� �Pp�������444��}P��a�����1��5�yjqk4cE������0���@��_��W(�NWܩ���W�QE1w�	vw����Ć�3�S���[���:���B��&���Q�>
�#�j�K���1�olmՀ�$����C���_����8c��m������QE�W�D"��MO��Z������D꣨�&�Y��`�J������Ӳ/Hͥ�Ӝ"�~G�����4p��42yꉬ[����1���@4r?�)�A�߿�@�
�RZZ
��| M��<M�v����:�#¢R9�7Q��WJ�����o���!/��4����iU@gam�.��X�E)B�������a�Ғc�9��3�ޛY��~�3ٳ����	���`�;����� Av��7XDv�Y���![�tj�A�V/}x����^4��^YY�����%�g�_��&�ڃ�K3p�_D�8E����)��oߌa�,�p^Ȅ���&2_f�]#�é���.+�D%b���}%��!���� TD@�7�h��77C;���� r����O�j����A�la9��q6x����X��� )̧������ Y=t5��㟙�qy����� �C�^s'H���	҃���;A�{�O�~�ͩ+4���TL+5ɮD������u�S�:nr��q�gP"Ҳ� �u���'������;G��Ӆ���������A'�җ�Y%��J�aH��鑑��l�O��o�[��Q�wHy�^����s�E��.�����g#K���e���kv+O�ͨS��%��-NǍ�7ުʫ4�?�:ihfXv��/����+ S���Ja/�E1KggaO//$g׾͕q���m�7G+P���O�`�d^=f7ȕk��j*��m�V��r������{���jjN|����ҵq�i��8	![���!s���q��뿋 q�5�=�rդ���M�eK;�a�mFbmc�G������[�!�d���rfQO�݌���vh�A���s��JK~rK$���&|6�ܿ���']���$V����<zD�"D���-�Vڪ�tއ�}�����\��S�
�~ų�]�l�J�H��R�P���7�sQ§���QY=*�\�uQq��,��O#'G쥧u�\p�B��1de	V{V_��\^�oOR!4.����$����*ռ�x�o`����]���ܗC�ev��Z�4���s��ϩ���jNn���ϱ��G�_|�1����_Qɮ40�Tk����]��uy���}����K��76�~5p�!eddx��q��{GI������c>�EQ|W���sr7;;9���"��;��=>��A�9�3�Ӭ��h�'���*y�F��S����-�KuBB���~-џU,��T�N4k���?4��]��w�Y�y7� kq_��������-_�Z�g���-11OW���[`2VSV6�v�N VTV��B����N�s�+8aa���R�S�_~Oq�����)�Lŷ�q�+����T8��H9�J���zf$��\��-nاPpIWnnA�W��3l�܃��8̎�'���b�s`ڞ���h|���UJ/�9�5����3L[�#����ɻ�N��:i����8�ȸ�gK]h��A'|`�G�Q��9��b`�K
j*�2N�{Lp�_�F�ϧ�d�,(Ł��6�����XV����!A}�.V]E��"�<�<�dlȮ�n�r����ñ�:a��*zj�����I%{�����/����"���LA\��!�ٹ9��_eo�XyWQm.W�c ��͓���!�s�������7��\B��}�&i���!�%��~��ص�� ����U@EJ�[� ��gu��u�MsdU	333hw��H|��'Y9:
.�`#�C�y3b�˙��0R�����O׹M�˖V��z]��R�\�x{�<�����E�_��Yڗ�7�c
���*�30�ǂ��.ͷ�K��օ})yzz"��X,nS�l#O���Z����ŝ��O�
��V\=|�-6�톼�Ω�ϛ񐾻�s{QL�N]�[�� �cX<7���E���ȇ�c��(�s a\,�-'Lp9����3�����$������āt���Ɣ4[�o��:��0���9k_�EY*��7���@ڲ��s�iNh��G��%�[��f���̀+���Ƀ�ۋ���Q��m��*0y�Z����p�����g�U� o/���|��K��Y(�����a�q�`pIE�3��̡�k�]D.���܃�Ϊ�F�g!x'�/���W�3�haE��?��OH����&R��}"�|��E��q0a������p��
�F>��f�=�b�S4��Aw
�FP͞���,y��s��Tf���B P�8Ҏߙ�Eyđ���S���B�g���v�_;�S3���V��?F�C�09��?O�<B �7 �&ir��nZ[���E�����쿧{AE�˓!��G3:(���+�ӗ
���-�ځ�0�򲺺����:��Q%����M�7������#��?^ܰ�/�5?C�Ȫ��r)�>��@y�ru���LFghЭ�F��H9�)~��g������˟Ù��נ��$O��SG�moL�������-�8�	p�.i����g\Y�ޏ���rs�_�a#W������P�1~ӕY��̝D/֞=pvN[i�`PD+b�B�țp.5��D���k�T	��p49��8E�N��>�$Μl��(����C ��%fAT����ߚ�V�q�_�?4��7�bT/�eE �!��E���W/��y�Iv�M�r��i[��==u�����2gf��;cy�d6������N�{>�]��Ŕ���ʉB��w�4��R$��F�涵?�]U'��St_B��N�'��	(J��a/1�8i�������)�'���d[�k�x�Df��:NŜWՏe]�|�?:3NLR�C�w��t3g����#^�׀�`=99�����1ʣө�J�����q�����"'&'��QeN'�&pBOܢ��|����'�FK�yZ�3[��FVX`�'&�l$/u��2C##)%�����p���gN<����㤧^:���Ύ.,j���A�����������X�[�,����lL�[�Ǥ�)����jAXV�[oI��d,-y�>c��Խ#@��'d����m�ւ���q?�=�c_�<��S���|�p�Okr�J����b��.�Kc>Z��W�uGBl����^��QNΓ2A�-
�K����<n�d#�'i̇p�HGC��*9�@�,���G�f�y$��B��ϗ��Ɯ�|�H��u���$���6���-�rH���#[��TV�WVV"���+ּ'2�P�3����ޞ�:���`�nTY7#%��<1������v�\�V����ܑj��g���5� Qg�毪ld<!���H�V�&99��} ��ƥ��"k��d�I'����#
�K9]�`m[�&א�ʉ�O�]U#�<(2\����BK]^b�'?	d�O*ߪ$����r�>՘�'o�bIu"����i���ͮ�+��.����!i�1~��~T��{2��#����Om&�3�3�)F��.9�
~*����}�r�kf�C
{N���pzf��_�;�|´"9Y������o{�8����G�{O��*�Aa��.�XXr���^[�	�\~���r��Q�;(�v־��+nܜ��<�ג�#��<(+[�`�K�˓?���y�ٹ�i�[�����(�S׀�����j�����ׯ_��(=�,��H��쐿B�^��~��f��M��K�&$N�.�6%FS2���,�ts+!��9�b;ѭ�$���$���ƯA�]Zy���'� �J��K���M$�Eu��7z*�7�n�]�K�FV�DI�h�5)2�����<	ڛ���8�0)��g�=zTT]�����h|�C�,��oc��R	_��W�v�ڧh�?	��➝�d$~'8��.�Z��z�S�n�H�#'�����(�J�4�Z�`��?��'rsϯ`;�S��4��19��u�'"z/^��ӪH�H�g��!��s�V�f�*{�\.�[3����C1j�������X���iE\h��GB6F��ƫr�U�%�ӝ�?<���^=l�}w��1ձ���C~~~q)���[���z�orEz�����9���r
�EGE�QS�����Şc)(*�e\���~a���!������?��
��Mer�<�>@�/�d�B��_H+����eG�EaA�Z���*TM�����z˔���!����B��C�PCL1~�HW�^j�����lw��~rB_O#�ww�+�UB����2���mp��9�rA紃��ږ�y��}}k��+�Н{��mY�D$�;�0p�/wcd����b;}���+��l���
���z!D2���S �������3EY�����4s�v�[���߮��Y`)O���v�{�;�.k�"d�~E��֊�	!��D�_��'USTE<b�n�+Ͱ �%�^]J�� y��9_w���ތ�e��w$$v
(��s�IX�3?;���"���'n��+�����!x"]�������9���;�;�@K�޼~���]�lY�G6����ծ�{v<�F�n�x���F{ɢR�����t�ș�v�8m�sS�p�D8i[�.�|��$���a5r����6	Mp	�Эo �������igS�z
�K��Q�� ���1.��0IqS�������S;�&��4ONR����~�O'o]@ �ڡ
��0�J���j.QD�N�U^>��2�����nn�]&�2g=q�����@g�i�`\�_�dQq�蚼H@�'Dl���N& ��_W~弻���#����-���B3���3Q�[���&؜��^3%J�p��B̃w��p�UB���]���Wt�c��8������|�d~>!�+mW> �B����$�wwߟ]V
�f���kp����S�,9��o�*�@J+z�5������_��x��@�����	p��c�� >�څ��p��؝����	����@ӭ�}�����I/+���������h�>�@�Va5�X{���!��=̎jz�5��I�$�@Y���+�ޕ�Iv}�1�z]P�z)��6��E�F�����_������\�Sq�w>B�|�\���X�K�[wMo!5����zV�<���+c_�.t���b&}Nr��#	�t�ƀy~W%E�(��k�2��W3�,;���L�#�OK/�Ͻ�~͘��o��}J���$��C�;}�����L$�`8�<e��3
#W�y������X	�d�^�ޚhO���Զ3�Zo��N#��^�C30V�2o�hkk�J���k�.<A�ଆ$bWzstr�v屑r���������|ŕ��-uuu��l���wn$:�I�J��=�nh�E�m�7(BB��gm��
z9���Q���Ao��|���7���/ǎX�$�yF������25	`/��㥃���5�:�|�~W�%e�d��z�\�J+ p?#�o}s�:+����Ԝ<�.0�	Bq�����K�Y�IcМ"O�D����5l^�C�s+�bD����@�U���v*�*V����ou��s"f�"����l 3גq��6�|
���)�|eee
͕��D^i���nD,�g��i�N�].�x_����΢�M���Ȼt� ����@�ۤ� ��Z���W��'K؁��h�Kj����2x��H�ʡ��
~�+���?_.�o^X~�����U�]���u'nZ����T���Y�}�?Ͼ��Wix �4<��E��V�mͷ{�~G�_I�g�Y���g1�Gg�%;�V=��P��"��)�Rύ|Pm�J�(�L�T�V��Y���:��{����O{�Pec�pjV?s4����M����ܕ;��ۺ�t*�i����3�b"c�q�Y��!}F���`��4�x�"��d��ٵ]���`�$+//���!L�=�0fg��@�D���#���xQ�ؐ#;��
�F�
�،~���5���~,�a0F߈9��zU;,J9m�,���>��2�-�����ŕ�@����Ϥ��L*ƃ�L��z����(��<k����?���u�p\��܌P��:)
�D��K�l�q[L�j���~MI;=u��D"�W2�4̌2W��:�DS}�6�qI6b�"���� ̸|�R�|s�l���ɀ!/z�K������
J��K��:Is`Z>��r����h��X���[PE�� 2�
r��x �ьhŰ�N���>a�J�#^P�!m��'�������G�J�G�(ө�����o3�l؀\� �6.�N�>�^깎'Vfq�U���H��Oƕ �Z�(�UR'�#�*�lO�`nR�����O�  ͚2�u�-d߫!����,A�B�izcw�<-b���̙��_�܍�*9�]D��o淜�tD��X��Ă�e�I�B�j���Bn�L������]#��yR�~�i��&��@1��&Ka��C4�3Fm������=��4e�������;�AD>��k��JI�nѮԸ�������݌Ù>��r�m��6ONNF���(G�l����pA��������#����&�������!�z���mm���Zq��Y�	M���=3K/{��\g�@S�z��@����bs�)'�K6��u\�3����<	f&����#�Y����7�O(��m��F�*�L�}=nrE�j%@e�yV>�ǙW�q4m�.;���h�p
��V�J	����OT E��h�:a>�J��q�gB��BRL�W__�i�#��An�6��GG�KU}�B,L�c��e?�qk:�v4�y��/˟>1yj��X��x;��[J�=��Kq��I.D���{���G�`�hŵܧ�{mO�8U��2Eʓ��i��d\�΄����fU���h��"n����u!t@'{���w��Ծ��w5���`���GoV�0!Z�$Ʃ�LN�v�b����p�� nP��rf�2(#�yz���݅��$J5�	g��]S0�@�S9>��CD�K*�F:>�D�U�
�h>۪k3���F�"p�������Ϻ��%���2m��rr�k��PSaQW%Y�0�\�s�_�ة�t�{���{���NJ1g����� �5$�0H�ڐ�LLL�E�ٓ��샔�t���m�P�F��g`����)x}�����=�"��_�����@�3(H)**JQ���.��Z� �E$Y�+g�V��3~S��u,C?nT��6;t�9�390qg��8��T��o����ˇ����t��e"���g%�����`wٔ��VJ��;��������b��h�P�����*�Bq�GF��jy�T��!9,;�fB YVv���y�؇�m<��'��Y?~����y���=��8EE8R{�Y�nk0�qFa���TT�؛���q��+MR��!�ֆhk���J���Tjo�æ)qK9�XfD)RǾ�?��H�b�-���ag#�I9���h��ڬ40���lB�G�W�M1�֟�w��#Վs�� =����oPCo�L7p��M����F[[C���A�F;7�7r
�VZ�lWUq��q ��t�~�`��#6�m(j@��?��Q���9��f]�C9{�&N�S�͍�fQ��-(�T @�/�q��i����R��st�{��us�x����g�����Z�ᵯ�r5�軿�t^ę?Iθr:�5�]6Kޜ#ݡW��[��*�S����T8��4]�]�mER�$k�i�ĲQ��qE̟r�2D�4}���.$�o����H2��ϐw�-mm���tR���T6
l���%k�v��#"�����J���H����Ut��z=�Y6��b����Q�]+�K�����|�C�ߏۤ`���.��P���SG�F�8�J㑝o>x�3W��t��ު���!�E��4��	��Vs:s��_)��+*�2IL�_�j9>:t��Ř�4''�Ժ^�RqO�q},C�ViB��?z=z�呃e�ѧF\i���(OÜ�8A�&UɜYڤ&~M���aN���uR�5�i�X$���܃?0��ʸ��~nnE3M=EDmM���T��DF����Y�/"�h��dHyä��s�4�h�"jt����u�>ߛxu/��NA�o7i�h;V��drݰ�_��Y�0��E��S��hR+(>K�E�C"�؄�%˯ �5�E�/OGc��^*Wz�~�&Tm`ϸ2-���m���]�wF�s��N�F���H��g|_s���t�U��&��x�~�-��}A�wa�~�,,�b��*��m�S��W1W5������f�h@g ���v[�KZ����%K-Sqal��2S�X�$%-�fF�.�v�fy�+qW�y�P���t7�`d8E��9֠-V�A�p�.�8,d;�Z�$
��u�\#j҇R5N���y��������sϳ<8w@���Q[>G������6ov���E���~�se���%\��|������O�=��n�>a��UTu��x�6��`���:��m����m\���ŀ�%��,�&V�a�����E�.;�J�@��}�w�{k�����>A':>�2��|]��I�ւ���`ᘉ�Z^,ճ�UW�ה<�sA�:�4�ϴuzQ����������G��^_�n�7�,����.�>��*l�l,7�?�Y?맄
���'�
GN,3�R���"�^@S#�4��9�4M��ܙ;z
�ddT��Y�m�ѡwwr�Ekp��FM�e)k,��!�<�&����P�h����V�ņk����$^$ͬ9�����n|��C�����Xw`��jy�1L�R��Xy�3�o�o��b��*�|H�N����fQ¯����/]e��b�����'��3�O}/p�T�`,�����oYZ��b(sޓ�0l1wf4�N�"�n�_ju�m��#*
y�������UQ�i��/����V��vږv�)񶁔y�r�	���m���~W8n�E�I	��,��.*�,�\,�E�ZAP��ϓⶈ�}T��L������ ������keA	��w8"L[�kk(c�v0�� U���z�e��wBN�6+ԕi�KSK�9��M�Pd �3y���� $�.��5����CJ\�D�N���<�4W�oBdS��BC.c�󤖾�J�C.Fj)�.��z�X��q�v__����
��ւ��*�B�������34h��w��=;i>q��u�<�ySS��$����4G����M-s�J\=A�}�m}�J�Ɵ#�M,��Ա�0R�A��U����T23�y!��!�N���k��E���*$@^�ܱ�>)/�BTm؏��%D@�fM�נ�Q����}0�������+������ZWܚ������
g>�f}�z��
6d����2�T_p[�\p ���N��)��R���� �v1h��<���*�4�f��l�������W�{�`tc.����j�]�8��RÁ���q<2c^�c�r���i���G�����U����D�y}j"lم�yN[�2���ozGc�]=�!E���%�X��-K��g�"gh[D�
����Z:�?=��Ɂ��ْ�/�9�T'{�oD�/�]ذ��5�n�;mzu�}��E`(A�t�biE)U)ڹ'�jE0��s��X�V
�u��ϻ��Xs��6d�]SZ�0��;,��4KK侠�b�dޯ$�50 `�8*s�ٿ ��i ;�O�EFln9�Hژ�p�B�ܝ�����5��i�3k����D_�M����(n��ɕ�g�t{������r��N�Baǃ��0	GO_@��YI��zjiy8���ت�_xE(v���e����<I╒�L���wdv9�󐪅�f��*^~��k�γ����u4F�"Jθ������13�U��G|�~��_��9�f�җ5<DZ�(?��I����x��0Ե��E��nK2�(�UR��ߧ��58w�C��;��HG���0��QpB����'�jყө��B�����wr�~���� �4�ۤ��[�uB�C�����{�eɚ�%U�TG�+�37xj��p�TVݪ1m�C?_c�A��=���эi+�O���y�&|�-bh�b̦]�I罾�X����@���@����~�P^�H�ᶁ����FY�p�YH	��c�X�#�;Pϋi!�JjY�;�{��kh���?���ײ�{L�G��Oq����g���[� QP_�+"�I��%���M%�y �0�c4\ޢ�@�������t��|��e�$j��� �V]���0�:����.�� j���0��e>'���h��ES	���T��%�-�Z��+�|l��rC��S�i�QP��{�!�n}��Սj��d��M��d���W���gn�@�"[���s͚ǿ7i�2�9L}1�1;"�L����j�:O{�<���Q���II�G���+9�:֑qGo'�/����
'��8r�$v9m�BG����.3冚�pE�u��ݳ��I�S��Zfھgjф5cb1��ߩ�PFRec֌���<V�p����uFD��n�|krX�-5\�a�\� �X2��r7Wd�(���,8��Z!@�� s'ӱ^*����:b�����x'��]B�l7��K��s�K�J�#�d�q���[��N+sF�t2j}ĒYw�gu9_��ؚi���㫜)��'��_h���	#�¦>�;q���?�*܊�ѩ����h�5)�˸�*��K�-�4���3:��;��|6��do���+T�<�ݏv�a'y���c��Ѓߺ�סnTL�*�r�� ���%�O�mYsje�8W�lV6�&.�R�땽��-��w��KL���w���w0�Y�>�2�h
 �,�fɦ��npi+��Q���ʪe��������BV��e�pr����9��'u��@�kd��o���� Չo�"�Χ� ������[I��i�&:�f&;f&�����Xj��1�Nі��@y�mn�q�uQYul�,��;i�n޽��c�L�������_9bÑg��|ṟv#<�?���[6�����4GY�`�D��	�;��P�"�U�2 �R:�k@*(�#�E?�_2��ob@l��nx���ŉ���n-�]�Mw3���`s�$��3�Yw����X`ى&�M�E F��F�T�</���ƟB I���mҎf�l;�Jk�s7�T��7ҍ�oY���pK��|(�,�Ǫ�e��
r�f����nym���aM�Q�D�{���I79��ʌ+���KǵX�聇`���lrRԆ�O&tU.��v�=��������sC)}S��Ѓ�0	�����/T#�D�c���22O�I7qB�S�! �Q��e�����t�n;��n���>u�1����=�|�<�8$ڻ�Q�/n�7u�2Ύ�My�V�E!�?�~�Z�'c��Fr���n��Zax07�4;|&[�#s�u7^+ȷ��7t��m��<_*c�8�j��n� n)�yM�0�?��7Is6���7-%���
�zAe\��-��EW�pf��ё��o�V���o�7�0�yW��f+Bs�ʼT_p�F�_��c���
����y�o� H�R0[�>�b�R��EǨsC$.a`.��*�ϙ_��P�4{�v2a@��ⶮ�G��)C�-0�O>�9E%@qq1Z��jx�N׭B���Nw��P���E���2f.t50 ��$�v��QB�����ƻ�xz'��D#����Bk��p��)]F��QU�q����iݘ���n��&�#�|�B��$����N84������P*H��d�6���P,3nw\��k����s冣��,��(��|�������|Z��Ƚ���o���d�/F�~Z�������3�0��{g�t�����0ċ�e�^�����t��%� �)jW^�<}· �˸}��Ћz�Y1S^.�`�+�����/)Rs������V�j�:���tD��t�hJ��=?$b&���D@���� �u)��2�7[�Ͽ�=��d��m�c;�@x�9WstQ�
�jJs��=�����C���Ug�b>p�:W |�$����@6��g�cB�h5�CB�T����-������~� ,�5 N|혃t�K�9��z��L�߰[#�u"��]�/\..=�*��eDpS+��Z��9�������gk,�'��w�����6�/�o�4J/�s<"ʮp�X�D��:�T��gw�M����:�3�d���j �9���9w0�+��r�D;Y+���JO8~����
N���A�7��p�jo�0g1U�j��˾އxn�ZB ����t���ZO"�u1o�����I�WVuZ
0��H����<����2	B�L��M��U!�X;p�o.�D��d�ۘ���k�B�����A���W�)��y�)7�!�y��0%��]
��;����@�W����<q�.���`cZ�0ckwV�u�y�x"��qoҁ�^�����H}7�獹;�a�N	�9��6 9$E�Tt�<�ޚ�{>�
���X0��;Br�6T���g�=co֨��� �j.��ۤk��lŞ�*���n��(q	n��xL��.�	�	�t�Ͼ�>[��&�ˈ��cwp�3�������E��~��w,6f��hl��5�����ξ��|&b�0=$t��~R}�~�w���}����z�o+e+�55�����-uv��W{�Թ�l��È0h��B���R��s̀��a����r�(�ߙ1u��u�1�T4cD��2��Z�c�2V��G��Hf�?���bym��nj�H�
��]i ����iR��U���Xϋ���Ձ̪b�\�Y��OY�ԧn���O=��òS%�kRQ��4���o�p�D���Ŀ��U]<����Siyّ@N
��#�y��X=�+n��'C��s}��J�l�߻oG�Zʌ�/�v='���t��u��.f��E	m���zI|`z�37�7��йJ�>��	��.)�ĨJ�B���*#��!�D;`슷ug�Cd�00�`7\���b�p=T؎��$r���:�jӝ�s�8�w�����}?��+~�UX�,Ĳ1u��\ᩐ7�;��ƥ��H%�n��4i�Z����~ȃ2�sw�?l���.���Fd��Ǿ�4Е�����0�~�9�8�<����$�3	(�� ~L�1�3G�3s��f44��L�uck�M�<��H�h��@8̊ü��#��'S@��`��L�S!M�S!��B�0�vKpx��B����g_��
��l��݊�;S����<�^��u�9~�)Iܜ��5�ʊ�V&u�>O.�pT!��qh��(����b���|�x@WË=�Vg�ʴb�~��2�:���0�N2�0�Ytn� _�B��T��0�mUR�vvx#�P���pm�pж�PM ;�.�~�.<d�w���?�rl�lM���0 <�J!���x���DW������
�gL�
w����ƧⲲ#�LC�o�Y]��px��loo�|��**p`��e�*�%~����x/�Dp|e�(�+iXk�ç>�d���*����֢�o���������&�]�V)�m�K���r���2��6���oP�/ d^ł|I8��Z�x�Too/~�'y7��YԼ��p�֚}U�lZ`���to��d�v�_XLۥ��v~fQ�_UY�	M"Y7��!�Uǜ۬�."rOB�C�Ⱦ��Z�!���:��~����1A�}+M�܇�&~ٴ�_����U�T�#�T����[�%ت�ȇUyZt}�?�Πi�3�-#��1~PzckSw\r*.��3��9�\
���İ��6l�L�`���"���G�m�����0n|����S]9����V���7�<6N+:9�ȧʹ;�����[I]A��4��/�*lS2y]���g��(@�{o���+1�C���νyZ��H�C�{���q��@E��'��G,pu<�{��T���ݸ�]z�.8����n["�Zض��������S�
�<<�L����p��W�������`��T����
�9c����E��J�-�6=�o�
\�ʁZ��%ϛ�͆^��EX9�Oh+���dZ��/�BZ�br��dе�#%"�q����<���^&J!���ɿ�ԑ�5ݝ��>��5�MK[;�6���XQu5'RUț��g�j/N/�rAc��Pg'�{�k@�1�F�ip(_�Jت�N�)�VZ�i#��0�M܏�{��aj���rB\;�u>�Յ�d��c�/�$��+F)Hq�D�Vz�q�Zu�4dO��"�7�z�x6���#1\_~y\@ȣ�z2s����j@�����\VnfF���h$�#��y&٤�%f��kG|@�V@������9���k��֕���7���!3�@�LQ��5ыӋS�#z�H��{�#~:B���3aży�PM��D�����.nY����Uo����2PF�n����n��v�ɍR����/�����E=Y��I�Y�/CO�*�f)K(cߗ6[(S�:���l��'K$aDC&{�ƾ��u�>���~^����=�v�y�����=���p+�K�8P0&����?p8I��#'g�r��m����������S�>���x$l�lؓ(R�3b��_:78�El���vy�1�&Jg��wS�-�A��r����Y�-=�~���v��|����5���#�Q�L�;�L�ѠrC�\�$�&��P����x�tH���s�h�;8X�Uy��ņ�F��n%+`���#��Gi�rU0�Γk��r���\y����o���"ڐp.��c��K��Y��SP޽�ӺJ��&���P��a����=6
�Y�O�ҡ��,��v��A�>gL?D��J��6v����mb��/��v���)��Mȗvݍo2�@����Q"=�[!r1H���������7C pЌ�+��f����g�}�X6�&�"�Q��Pdz��a��K�h���#?�_�xh�[Ѧ�B�׈������˼_��~T.\>/m�R>����{��UO�8�1���V7M�Cz�F����s� ,H����&v�k���7�7��Nw�qw߇�u�G͛�#���I�"Wt�$���R $|��:�Tzvw��&d/:c���u�^[�c�{myR)��ģc؉\=��_�6�)�޽o.З��K޸�ImJ�\�V4b��/M|��=Cp�#�#�o��g���2���wT"	��89X����[��Vhڧ�T�TXw�T�o�����.����')��;�@����+�H|�	p�D�
l�
l3z<q�����Rҽ���2D�� ��V��O�=�5S̝R� Q��-�ޫK�63��f�1����^@R&��g����OM�����R�9�[�I3�\���)bJ�&��>�� R#%��T�8d����L�@�����o�X�w���L�E�HH��gE��Զ�:l��0bcb���3\
��@`��u]g_��3:U��iں��,�[�h/��_Hwd�~@_�Up�T��j��wi�m�<�2�i�G��Z0ń������!^�]6�N%e����8ڣl�@��*��TӨ๣�N��d�r/�-O�H	�ЩO�}<��� �|�S�����D�q��ڭ������55�N��i��m�Y��aHf��4HH��6Ҝ�w��D?$d�lz�ۍI8M���j~2������k�.�"����JöO�/��p�� �m�t�Ɯ�X�g�#����y�9������%H�s�%�b�c'T�] �Nwt��Ap��n4]�T�b�#~1�vk��T�G������Y0�#��̨s������Ndy���`��m�[�Ȇ��k`(S��k��DHBv���*?��v7̡DWg�Ǫ�0l��?�D���݀���.St�'�K0j�jLR�	�������3����R�2H��Uh��z�� �Y�R�����3�uKJA�N}���z2��Mvǜ�WɃQ�}`BŲ�@ѧ������1�%~�O/2�ȑݛ���χv������tF�,V聆N3XS��������e�S1	M$���� >��3�%2j�������~*���HZf�;�NF&~��n�7���W�#w��5i�ſ���]ʙ��x����=X:�΀�'Mw��H�1��m7ġmr�D+���v��k�6�l�������:���ƾ�7u����p�ǐ�`��{f�2S��W��o�m���N6�c�OXAC#Fk˓�/��g5~��vR�'bD:,�\�R��%u�\�ᝉT�L�������ҫ�	��Z_���-:s�M��Y+og��1��=v�b���S:dӛ�����o�'`}����_��_�j
v�W��څ5���~�5w�����><y��ykĝn�)%.K0�<s�y�4M׮5Al�|�qv}4���Y�|�@���	��1�p2"�}&���X�w<��r^������\mfw�cg;�܀�?e�\%�0�a�NףAΖ��+9�;\(\�d��카0mk����H&��8���M��`���4	���r�X ����x�ٶn�8����e���_Z�R�'�	>	g���e���R+&/�����C���3ܯ�cTQʏ�D�kK~���É~
���Sq�v�8�	}���;OKW^n�@4�ia�ux[3�o_R�������\	�[�`�PRk_�v[%u�������0�d������z�x�%�������
�$r��
/	*v��+|Ǥ��oW��u�5E:w�ڑ���3B%qJ|�E�P���a:�r_��:�ej~���S�?� �r%v����Y��D2ymQ�q��f�R�x�ل}����=�3c��i��
�7����M��]>�T��X-��!��ۍ�0���+t�$4 �{��n���Zٷ^��E��8�S�1���GB-D�ٸ*c�R("��������mA��R�{��G)b�D��c���|��u��h�Yg�b���R����GچJO]����b�G�|uw����	�����N�����Q����._p�a\��v�FԊ�;m:U��m�5h_8J9&@\��b�
f��#	�c{w/+^mn@��L�Ë��Ow�Mu�c�s�]���!�I+��_\��'�2?���rF�p���C�
,y�'��oS�f�h���<UjW=��E��L<�	 ~��:���T�E
3����Q��\�}(GB�P�d��X�3��!B�;�����
ǃ�Mʑ�Վ�f���m����o�� chnf��IͤԶ!��Pxr�I��(���6�	�\Q�������.�FH\��T
��m��NQ�;_:҇H:eԦ���÷��'�Tp�OUkf�` �t)��� �� V�E�@�(�͆OaF$�н׷))akx�������ԛ��Ԩ�.���R�7���Y#M# ��:ɜ�տ�4S�۩Q�1��՘g�R��g2B+p��>��)��{k��ڪn�m+!P1U�awO��ٯ��7?��=��f3��XK�$� ٝ�>��I���ox��~^�X���.�]�&'=�{wͭ�;E#�� �����O쀠:��p���6���j0c(a`|����EgE;�u̦�ef߭��U/̬��4�5ض�哝?�4�����tS?�m�C�o9�Jh�LMy��M\Iy��8�{k�+�!V��蔊��)ͯ��6!u Yϔ�>
�4���cXX��7�g�p�d���9��*�m���w=����'�Ab�'�:Okh�6n����p��<�mյB��M1�b��lIz�u���`}�{�+�\�~�E��� �Q���36�I�Iķ'�qH^���$Z�27�'x����Q���T<��5�X >Tj���d�w�h0�N̉�=w��#�皎�%�;Z�P�
�xK���O;\��i!m���?v�����&��e�ªٴ�ݴ3�����i*M�2	�r5�����=Iȼ��ёI���?����1�~�,��B�K�Fa]�-���$�Y�Mx��0�y?��nZ�Κg�Z��#���z므r�f�410��}~n����}�'L3� 6>O��.d1j "��)5���U�D���h�]�G�%��g��ە�G[Z�W������:�?��28�ݛh�"qB����_��͗�E8��k�mw�"��e��]��@���D�ؼ��6ڞ|MRvƷrI)���V�8�`�k�)%���.k���^�; |/n؝���е�������0n(�gh��Ǝ�[�NJ)=�#{�Ǹh��j������Q;L8��:��c�*e�)^@����Ej3c��A{B��4�oy��~l��:/{oS9u�u��׊`�+�{��Ԝ �Ƙqї��@T��OvHF~��1>��w�`�����~>�W^�=�.A:��.DR6|i�]��ʤf�F���ϭ��#6V�cK�C. �u�{��r!^9Q&�:����P���}�����k͓XW'�L�Ee <�[�R��D�΢�<�0�P��,,�h[��� t`�X�"{��8�R��Ҩ��F�>>̛��i ���i�Hi�m�AL�\���z�/���7?~�$}��}�]������Y�т?ql�rf�I�'�a�����G��Ѩ})�a�X��i�&�'��78����=���
�F����F{��O��qL�䚿n��s=$�� ��,�}�O|kKBgy�
+���Y��b�܀�hWL5�0��Y�ߨC<�����!��%!"J�?=���m���SH9��b�n���'7b��m�������A�Ƹ��^%,Z�6��4�4T4�y�v�e$�w���:xm���Ҩ��EN�?�[zR4����v�*�1��U)e��hsr�:�PD���~z�?���A�L:�7�ق�s���6�����f���TC���^7�}i= /*9eP���q[8�(i�4�u>�5Iv�ٚd��ʜ��t� ���#	�,��#k�a�ܣ���k����l��ׂ`�	��+���T�io���+å�.��3��6��z!x�C�
B�"\�W%fr���Kx�Q�'��i�u��x��z���UYb����M��t��L���ib�wT\R���ֹ����F="W��͕k���Í(�����&�4!�<��#��l��f�5����7׏�����f�6%�+�� -�ع�eR���P��@�G�F/:�-��̷o�n\����~�4cg���F}����à|P��H��I�����+aG��:��� �2�	Lzb���m����(҃����
�A�5�A�q��?�e�7��~:7+��(Gh��AIhcM��<�'$O�xEՌ#�"�T�ڜ(.Jd��$�|�:��U��+>+\=?�Y1	�R���Ǻ\������U�h@�pa�{
��5ר�d �6(��|�Q��5 ���_^@��R8WOk��mjz�Goi:��Z�݆��vg;����@]`���̮ɏ�~!�]�?W�vs(�Aè��m�u�Q�.�g�0yAj�6y7{AEM-���;l�4@ L$Hv��'�6�H���3�B��<GB,H#/.���kGB�ɘ�k�k:tJ���U���뇶�S-�+�d�=D�*4++-<�v�^�j��k9���gp	@P#Q�$~>,��?�{�u��D�	}%��O�'.}� �{��9Yl©����c�+19�ϡ�Z�>�:�^�ư���¯�I,#�/��|Jy4�	ہwqLT�]��T��WY���W�E�/"�y<��z���~���Hw���0�ܼ�� ,�U�ٿ~MMz�\O�6��[��W&�SxW6���� `�G������ڑ��b���\3�U��X��-f�au��P^���h���(�@o��]������Y�nj�F��f�C5mBT!H�� -�,�v��$��]��
���z�e�3Hj,���n�))�����/��E�\]�A̬��Ö�Q[y��=Õ�K�/��M�q�C���c<�w�:���^[Q��l��^��?u���ݴ�R�ɪ�&�ׁ�^�K��wٱ_9:��[Q:��(�m�KM��I�7H��'Y��C�
�A�Z�� �"[i�4�m��LT?�)7t=\�g�*�yH�;>�T# Kͷ�O��������:���^hF_"����d�ڢgo5��aL��S�HB�a�0->�jI��}����{c�D��T���|I����*}���-.�^���L�T��C?7�����O�veM��鉮�1	�Ž�l�튱����/S "��y.�~��1���v�.�S0ٻ��B����F�u�4�Ԍ
���3˟�O4@���
lۓHR�ъA��S�'�G-�kE����6`Jdg���ԶLao���ך�0�%A� D��*m���itn��kF'�;@�Qc�8{���z��m�U��):�,_�K�X�]�����!36�F�v�{�5����n��\C#�82��qn#ړ@����f:W�q�Kv��D[��bӛ�ׯo����q��9�~g2ɢ�<:�m}l0Iﰮ�4�HǵJ�����3d�t�_� ��|�l����t�Y ��o���A����9��R��Ql�U�t]��ѫM��V�VMz���c��a0�H��BU���He���
�%�{y���p�(K`�����$_S��/����&������Y/bw��F��{
�����ը���Ro~J�͘��~pu+m�|�5QK������@~��W�5�>�h��j�)�jWB��x�w`2�%%��YVF��
���s�K&Y��|�m�ػ\���s��SjZ
�{��{�#k��#Ǭ��^��z��Ð�R��m�X�e�:���lBu&�f�q�T$MR���dl<����5��|�J0����nr`*�O����p�[`��v���B(�[u����s8D���g��NEQv��h��ڇ�q~�(t�������rr��;�'��&�]*��]b��I�g���&��)Sǫq��yk>7�|���j�����m��Lv�sy����-��Hg�I��ZT��A2�^��u���F阜��8v+�_B�o�~�u��'��Ҟ��#��d���[O����S~q:U��*0M��tX�M�[�hM.����<sϠ���4;UuvB6��CM(f�T�ʃ�2������6ss��T����!���Mh�5��ѭR�
H�Z��=�3��Z����{�Q�b�L3�6PE?J�wt�(�i�9b�K1]x�(�Gf�}����C@��^��9��x�[*m�|�h�i��lO�#mV#h�ޱܻlݦ�[^.|���Yi~y	��8�;P�RV�wZ�0�^0�jz�:� )�k�I�J�&�;v0nl]��]��p�B܎�u�L�w���W��Lռ5N}�}�/����S0J7U�Zo��٪E�S	}�9JV�H�ωR�~3�#L�W�r��	�}#���IƶcG�d����#&��B�@ƾ�K�W"�����.���X�����S�Cu�۩��A�[�gwj36W@���):fȪ���T@B"\�
��IX%T�h�D<V=/S�a�J�^x"����2V^}���VO�l�k�v뷕Fe"��u���������ָ��&���U� �*+z�9*�־�J$��Mg��Sst��<���A��F��}�?8w{I
���٭�|�@�$m�E�I̦�`:f�:�5$�@P�*���=ڧj��v�XJw�0{:�����?���_i]�4	��m�R��M�k�c�{�kQsjOV�B�?��L�'JL}F�w���ϯ~���p��L�(�=�j�(�6zŷ��[f��P�3���!�؜-�� �+�j�xJ��:oL3�g���v2c%��tO��Ӗ���4J���՛?r�o�1.��~�I S����_z������*a�_ص��e�#�K�b�=�_�r�9=?�Y�,a�v��vSit$���o�
2`1G��`���"���T�V��/,`�h��kv�6��� �맃�N+�{룷�uk.k�l!~*�.��h%�{��f�`��^[({��Cۓ��X�m̨�S������ԭ���V��E!qshh������`����h�I���b�u�/� ���#��>��I���2ִi�I)
Vpw`��Th�&6ME�;��G���/ߥg`���r�2'S��8���~g"*�_A��ϙVȌ�ϧ��Q]�0*Kn�('�g��lp��?��E�Cη��buW���/z�m�l��GJ�śh�"��P�� ب��i��P֘�*CF�{J'`�T� ��{�B#w&�c/�Ri�����b[ƶ��"�	��q���H��(���y`eQ�(GW�j%і�]�S	�f����\+݈��O��y�l5�e+�e%4��/�ĺ��&ϣ���N�I�&��&y�V�pk����ҏ���s�l�ۗ�*�ZG�81����-zX�:;�����ؚ'u�qп�o�L�FRv�Г�]��S��7�:�T�*ޢ6|��=��]1�����z1qu\ϐ�9�&z	�B�z�7�+�J�,Xk�ݕ�X���^j�>T�&�On�rB�mc=�����ы?�={A/�"�
xl6~���;q����1yĘ�i�(�f��?�vw��1^�Ѱ���x�$c��/S�JJ?Ȍ}�{A�xxz'$��w�~���]H��e�����e��6!������D[� ��V�Q@_�@c7�?�a��<�1�gΓ�,��F�*/���{V�5n[��W���Y&�cuf5{h�>8`�V{yY��h&U?gpE�K;�����`�Fڎl��-��觉���p*��;M���D�ˊ��7�MZ{�I+��E��1�� Q�Uѧ����7Ƃ�Ǥ������]s��}��Q\�܉��S-��Dq,�����2vw�\������F�����i�?FJ�g�3�]���2��w��ܲ��M���ں�k��������0��܆x�yo���Xy��{3����e���=���3Jێ��ti/󜘞_���N���?=?�)����@��NSg}�B�r�7�T�P��]j����[�3eV�;$[Ĕ�|U�َ�I��f~��l����]{AƩ/�,�f�*���	O�`=]5 ��cv{��Ġ�3?"0Px�>6`���2n� �q���'��tg��[M���7k�	�|j<ȓڬ��P�P�������Ȏ�H�4�vw�|��r��֛���jD��R���ϟ�V� %y���� |^�����\lM������/_|d=V�3�����g�V�V�[����e���_�qH��
��pͬF��z���:��M�PAr~bS���/
'7:r�i/��HN5M���XoG�iy	��-���B����"�]�V�@v�T���-V{��IYѭ"O�/�,)�b%Z����y/ɼ�͘+����F�R'�������F�nr:�ԥ���旊��u�����C���Wu��p����:ۖ�w\f�#7��Jb�x<E;�'�wr�F������I_:�r�t��HΫ�7)#kmZ;��>}��b�����]a��Oц4TkN��>h�?�*>F�xz(?ODt���Gd�OU��1����Y��WO3{����|�U�uM�}�4{��K�_8/q�|����ϵwhv����ٜ��"�H���s�L��m���O�On�޳ek��rp�o�ݲ��N��A�s��U{��t4~��o���"Q[�2�0����NG�̽��X��M;JC�_u��� a��G3z忭��¤��#���e���u�_:
��X�7��E=�Ͽ��f���vO��a�L�NL��o����}a�TZї��ηi��LRrZ	Ur��a���<�������V�]#���fd.A,�~�r/y����A���|��P%ɪ��9�"�4g�^eu䛟��<�J܃|I@ٰ
�Z��:4O_����	��e?�.��C0:�ȷ��벢�6��3S?��Xy�/�;�ټ���q[SP��d�S��/�w����e;�#�W�����=ZT"�t�>9�[|����9[Bo��RQ`�+�I	���b��֮�晳��Ri��/Il���#��,�~�����q�H�����X���	{M$��<��ZN{�b�ϛ��򒚤�;>�ݫ�Jp6��fOӯ]�YK�D�s��<���H����o㴣����������|�M�o�Rn}S�A��K�*�3�����ۢ�z����J.mg���v��f�ds��f����a�w��=��:�����f�Z��bx��a�oJ�����l�H���眓�X��zy��0����|>�+��O5�;����Kw����THxq�.�̰YFX��ŭz���=��������7Q�v�QF�����%�f�])�\9.�;_��Z��:Ŝ�j�r~�����Z�cj��x���A8���Sn�*�m��Z�;�K�ּ�������Ծ����r���E��xŐ��f�s�/3�aߖ_�I�J�	�e�� DݓS���>�͸� 5̆�z�z���o�����FT�Cf����)
�8�8n�O_|�/��=��(�/��#�_��������&�ݎ�2U:%��Cs�(j�*G~]�wq'D1�""¿�_�$/���J��E�Z�b��~'HT�lG�jӐ�=O�b��	��Z�8����׫�LR���VuU��H�A2�M�b���Fᆿ��"�}����-�6�~�b�`f����Js�}՛��6_"؎��X<���>?y�&"�{E�����+�����Y3���VS������Άt�j�[\��P��Ȣ^�����,Di	�oS�Y�^�}?ѽ�J��-,��O�{�A{�z��(�7yb�?9������U�$A�X[{�L�~GX���"�DI�)�E}�af}��
 �]�|ļsӻhCmΒ$d��M"9�R6��!}��i�)u�S���P���_��b1�g�`���q@7H"��n�]Z�>�`,�)$�X�y�ƽK��E�~҃�^�u�+��K�G0t�HD�����[�
v��`�T������X"�s�E��+9���;�j� ���@�~X*̞e�ڲ�V3���r���"&d��5�R	���;7K �𗮎����<S\.�ٶu���W*sD���T�z�DIuO�X`m���.�8�
��#�����5��O�9��f4%6�=H�v�]l5p^�'�,j�_3��n8� 
ͦ�?���q��\��^�ߔ���	͊g��!wR�3A�n5��/���]������EP�n6@�BQ�}#S\�0�Eb�����ѧ\�B̹���_\��֍�N���_s�(r����^��e�!v���<���p��2R�ϥ���ې������M�-.�ѧ22�o)�R0��s{�IӇ�^U�G ��y�	Ue����<S��oat1�~��SK׮�|�sG��őg�!,������˄��Hw%��_v�Z������J]D�I���j���¡�	8R�*m�)��t}B��R�x��_�.�R��	N;�ѯ�H�u���i��U��j�x����ń>�nT-/���44L�c�2�)&S	�{cݯ��=m`���@�B�K�Z���NX��B�v�qi}�Qv�7�<μ��"���\��u����J�M(�O�	9f�]C<������H՘vҺs�N�L�'�k0�5e�oǳu}˞-r*P_�����kDw�R��F��"A��GvZ���FᮯJ�xPn���K�O�e�Bк��]�˛d9Sek�x��o�wۅ���s�-�ɜ�)F^8�Ѝ}:�%��10m.	F�ͷ��<�Eb�@B�������;���X����ؽ�#��_�s�T�~���L
��=J��I~c����UǆU��v�J��J��={��r:��!ۊ�E���mB������ZW��<hV�،�u���z!���bc��������k�i=(w�K���"��QQ.���V������+�bx8y,rr��!��Z` ���G�ЁC�?�J��^�JD,� ��B��lM��$y�e���8�c�.
�����P!��)G� :=�a��}u�e�P�Ÿ�6�������^����}�Y|�k�*4��k����]r�7o�fS�i�I	��}Nσ��]��<+�
��0j%�[z���u���r��%5 �$�]�l�I{ej�x
Y��w�f�"^���h��2�C xֺb��Ż��"o���ߠ*�k��?tΟ0�Go�J ��[\HA���i���4
�-[�D��W?�M��i1����Y�}�
g��s����f{���KҪ'y	�ϗ\��;Wh�e��J4a��A"�2�t7jELy�����,>[�� ӼS�l��rd���ʙP��F�L䌆��=����䙍��+�������F��A�%�%�M=�:�R���av��o�{o�/.���s˄Y8^�:r>�P��vX*n'�T�v����l�={��������������L#�]��b��rE������� ��Hحu�ð)���D�uBӯ�w�rxfww[�(��q[�w��t�Z�yi}̃+�i�zdξ=�ɂi(ϣ�6L���Լ��e��@ Nr�N���h������j�(��UcL'�� �3o��b�v�=~������q��i�#ݫr~���C�Ѓ�>9��8*�ܮ~>g'EW��#�{Uj�Gd�� ?�]_��� ;�V�����l�!�T���JB���5Ӡy���{��T�%��Q���4?w����DiT���w�o*���s���={�.r��qI����f��r�F'x=A�}0�oa�t#��h-W��{��&�@J�����Rˎ]�n,b��������3'�E�=,l�)�C�Z&8n~X�<���% '��?�O�f���ųncy�rr�� ���q�����,���\�t�Ӎ� |��7�i�5�t�Σ�sZb勔j�\�]�y��g� �8S"�.�Y9�:!Զ[�r�o3b$b1ۗ>�r[���F\JZҲ�����i�Xȇ��jLV���Ɇ���	8E�����fůʯ{3�0��Pv �&NE)�>��tNtK��F��V1I�.��r;G��{#��aS�$��k��	�y��X��Dk�â�c�P���H��ZK���xut�Q���;��_��*]7��__�?e��|m�$GD�o&����
��i�S7
?X�
e�<p(��W�_�Q�/�d���3!,��Ig,nh������DFjGl7�	��oX��f&�H�DI��oۦ]>4ג�6.�_[��~�(X��/�p��l��vw��q�"3�C|�X�H�����Q|�##��F!gf)Ϟ�\�Q�e�����h��v\(�s�-�S}=���ǅ�.~(�r��"`v�|�A�NN�⏏'��_���2����UE�/^�_jt`�2��Ga��v7�W ��'�]{�����j~;)R���rǰw~�fJ-��a����uY{���w�LNP�5�k�;;g����ԃ��#�}��/��t�m��ܤ��|���2
���c��y#�W�p;�l�����޽K�t E��{����45?��D�����d�z�8��>4�m���/ҧ/ہ{h��E�Q0�F�r���op56V����6s�N沰Q6	�|�#IKU���g����r�MJ�X���� ne��/�K$� ^����t���L,`{���3>��8-���:j�1BQ���������~���"(M��z"�2X������N����1�j��A3?����,(
$�?f���VW�"2	���f>>�sgs֬Ag	r_s_n<_9��#�"p�E�P�`� ��ip��	�R�ŋ��7j'���˫���G��>>����N��4�zl�:����I�Z|  å6�NU<��}&f��ɖO�R)T��u��������"K�s����/S�{��q)r��Q}^3t{N:��/����L���~��E���ğ����ݒ��>x���8��e"E������+�o��g��2�?��i��B��w�Y�A.ǣ��L���r�+a�
0�lb�|�%P=K��E]���EB�^��`bq�e�ݾ�x��ZGt�=KE����G�(ח��Y��C���3� �<ˊ��N��٩��3M|d�6��~��^:�7"S�G��[E䡕e*�k/��%��;�׆B��u�v����?K��ֈOC��Bq�����g�~"y��-��Ew���p2m���y	\k�5У�w��+l\��Fn�[	�ʶ���
<#盥�kb!�4�b]�T�U�u��x�[֧ϻƋ)S���Qݡ����,�Z���*���p���C����c?6�����I$g葿ZH�w�-�)6�#aa���|~�ߍ����y�R)���&,g�2�G
&1���)�D}~����0C7R\/o���D��ERzQd��	��e�~��I�����g�w%s�=5Bf:�0�J*z�d����>n�㵿Ӯ `����0Z��TsK��ӄ[
0�MS&U�z���
,q�D|C7tkvP�>{x���8�ZI\$,�g�L܂����� ԣI�%wp<����`�X�螋���$�E@=j��Ȣ#��oE���&M��.��-5��O��Se������?돃n�ll�7�Wu��~���ˢ�d"YKC�O��Kx5��H��tm��ӮqȾ���5���1��9�]�y!��I^�1�ySa�1��t�U���۳c�����1�n|�y��<܍ɨ�/[������˶����&f<hM��3��č�0�A刷Q2%u>� Ѐ�Hn���.��cf5���(�4 �w�!'$J0n��#��@3fi^Qі��l��P�p��S��A0�L�Fd�3�>��#W\56zmݸž!��tJ�r���H*4��E�h��x)��<s�����ܝ����do]2��Q�}�ǲz�T���CVP� 6�ySc���q^m$�!j$��1wX�7P���*[y�}�n���;�"�`�bբ�޻	��؎w�2t��y�R���JטDB����QWoj��~U�N���bT�9Q�f��{�l�bӫ�Ս"Y�v!I�4��^�q~����[��U]������"Xe��N��7��aJ��*h�n~�F�(��s,	���5,is!��]�<�������y/6��N�����(W����0����bҵk>��i�%ի��G
1�hܕ�=�ͭ����	�4�B���i	��;)�_R���q�HҨGH���5x�z,	dfG�@ZZ�al�a����#sroS�G�GT�H&�Q=���Wj�ު\���UĠ$�Y}K̬����P�����M����=޵���*���Q��u0�,NS�{��b�L9��o|<Gk�Dk&���y	�~5M��]�1'�`J���p����&Y�����k�L�t��JI���3��OAD��w����T:kMBS����L�ZӁ�t��Q�X���M�Q�>EBg��ܺ-�� �		���94���a�<�|^=���Kw�Og�b\-kū꽾&��X7`�3��i1��іm�+��d�(�w���A��DɅ�wB�ǢF�W˾��T�x})�DN,�G�y�-��= �E�@
ī)�ZJ�f:� �1�6 ���_\f�h��Lf��&$>CdִӖ, !w�$k�d�&����-�!$��t�W��%�󐋟A#˝��3 1���Ȣ%�·$�=�X���J���ɽ���B��0���������¨n���޻��֯'H���?�hh�Z�3�����������x��!����9�c���CX�$��	�{�D���b�2��H��q}<_!b ��p}׸=y�-t%$$D|���g��ᡞJ�����pZT���g��Y����͌ݖ$$I7�"�>br)/��z�O��k��%y��(6�HA+�t�c�;s�$�-usC�ޘpeȅ1s�+M{�h��h
�z� T <���훼�N��s*x�0j��DQ�vU���s���.�Ua�T[�o��
���	 ���lj�1���.n��"���Kt>K�ۺϦw�|'%��ܟ�)�Urb�����q���_]3��a~�А��qCA�X�Ri�=�5E�۱nh
�(��e�������`�1���#����!w�1��x ��L&E6�!��|͋y`m�tg��j��DJ�|pOu��0�^����q:��X��=��3 U�;'�[y�)Az�;4�����ڱ���eK&��G��g�'Y!�=�ԑ[�UB��� 3�*s��gN(V��W{{�C#�S}����
���:xЃV؃]��E�a�#�X`	�����5V�_��������t�e�^�\{�#���xș)e�WW��36���U�SL�����D���͙Xx��`9��Y���?������-	��)0n�m3_���n��ꥯ�w���L=�(u�.|�
C�-�=��L��ڍ�rL�1$Tl.�������y&c#Ƀ�4sN/�+��@�R*cu���,=��9�4sz�l�N&�X��˦;���8��Xj�#��UQπW��h������L�8		*�X�W6�t(����0b�X�,�zf<���)�_�1wu��9��(1��(�%*�=沯Z�"�<����5g'�1hz��i�1�'O����D��5#��)>�����#�@#4�$��	�͈��c��s$|��d��Q@�Ni�E"��]�?�yAj�旂3��h^X����OK*�t֏��i,�0@m�B��q�@��1b?����y+��}���و翵p�<���|��d��=fQh0g7B�US��� �zV\����'aRB���P�'U����?Z�̺Y�&K�k�#�l��)=Z`�#߿�ߧ�6��26.+uQ�l#���<y׸�_�7�5訣�V�:W���XHmjR��g "�9�6ײ +��v�����]�FK��/z�G9����]~�&��+М^;f�)t�-���tR�a�uY��ꡡm����/���~�t�����TӋF�5�ͿDy�����qf况[		E�Z-�Ӈ�\���QF`����r,"z�b���0a#��t��^�{���`��c��I���2;D�~@��fi����/7�͖�_'je@.�A�0�<�L��̹sg����{�& 
&Ix_�x�F#�",���:������SF�mvDy�<,�'(��������W���/]�1�����Ud��7��c�����9߲X�}9(����*��
a�|<©�83�`L��oE�T��=��{�}I��w|\�6p�O�:������U���������S��� �Q���.����dW���]]�[�*���;���ޤ-��=����S$.�p57��Yt��mwO�U;/Y�_I�T�L,`p)"#�/(ۑܕ�Z176�{\M��\"1���L:U�?�'k�C-��>=$�+~���v���*wM�35B��]���󌋰�d�ֵb�!��%\��υ:㢒�|�u\������<��Jz�N�Nt������`\TF'�ݪ�������>�Ee�j�[0N:8�Y����b\��q�ӳ� ��ڱr��%�\����?�yD��NN%�7�k�:Ӯpx�.��Z|���ۓ�EB�2�GK��ݓFOA��dN����4z�J��ْ������o<���A�B/&��,�aEB!�0��m���.����/�QbhhT5�qC�}m��;m�aC���MԄ�5 <�m��w��N�oU�O��`Q[0%�6��&x�)���K�l+�<e�ڂ)��!��1��^�)^_�3����L��S��/���,h�4�)ʸ�%Ꞇ{�����������Th�Z��?ѯQ����z�ߘwh5�\�ܓ��s���D��nH���>��ziM�s��q��,�ҥ�Ax�����nlE��c{��{�_9�dH)�,���L�-��'\��]P4!HG�E�%]�&��n�M�$���F�stvD�W�s�	�;)'|�j�d���h�)P)h�C��;t���}y�M��9�"�)���3o�A�2�o�3���5�T�H�j۽X��TM�X��"��	n��!e�����l�p�1S��2b�ԅٙ�}���9��svR��q�-���FiR���Z~�	3m�l�a�Vm��	�`\���lV<��B�D���#t1�ty|�����u�/vv���bV���g�r�۞�tt��y�-�hQʡ����;W��ZFFz�亳"��b_=��_;_�3H�n��KK+�*C:�q��I+���^��Ԁ_�>��%��jbn��	*Ј�^�o[9_8@&ʦ6�*[�^	�Ill����\O�[�$ ��{)Y�o݇�X��ԉ0�ԔoY�Q�Ua�	>�~7��-�{_�/7TG}�
�r�~���"ˑ��~��k9���_B*0�9ـ� ��V�ik�|&Ωy��|��s~~z��h=䴰ԨnpN���2r+z�z�c:_���<E|l��DCJ�7YᄄL{����� \��׌q�vg��Fg c�N��Xi�����􀻡���&}�c�:'�E�2 ��a��ɪ<2��x�
D���x��V~�
��R{��hgO�7�#�n(*��T��'[m,fQ8��?.[��Sd����q����A?���H��,�:嫅�	>�	���E��a��#ۗ;���,�wᵎ�N&U�	�\O/b�|F���J�ʿ����1deJ�dU/�%b���j�q�!4��R�5��(���J'�UMy-���=3�:�zc`N���!���x!e��8/cX����
��5>z�M��/F��>tS�֚\P&�R����=��&�����w���ϮPܧ�-�-�z����3���gHpx�z�/�h��X
�I�jq�*�{+c-5��o��7�b�r��S@#��3����Bo��?f�b��lF�!��@/�T��Yn��kƱy�ut4YYIg\{O�*>V�Z���}����6����-z�L�X	�0��)�������;)]�Vl����|�� Ӑ�䭾���fXdG��}nl����7�
��V'Q_k�1̢�%���Vt4���SUݢ��w�t��٥���d���>�'��1����8�E՟�Gi^K��y�-½����O�zg�V!�~����q�Fq�� 6���֛B��㖢M��(��Td�,�-JE܈�T�컬ck���2���.KʚYÈ�2ٳo�{�����}~��y����9�q��<�׳�%�Pp`l������˾j0�q�
|t��J��)y6lΰ�W��﯐��7��Y5���i�Lɻ��+�`�}���w���/!�ڻ�WM����؟=80F�@���^�
Xy2@&�~<y��;�=0΂�T� �<s>l�/�e� I��>�%8��;[����9����IH�9z�k�h�����S����4��+r����`,�����4lnbB�R>��x��
�MM>W�*q7y�B��Ws�*׋Ϛ�.'{��lKgK����A��ݶ<R'�'�s���bn���%�x:���r�� ���?-IW�$�*2 ,<��?������.�|��M���v�$��!�q�|�j��'�<@u}��N�]!�8y�����b�]R�]ѯf��pMN����"­��I5������`��KS�k����d��$��wvB�%\PŞ�9��� FC�z�myJㄉc�U0�=�u/V���"SY1jF��)@�'c��x��+��y�vL|��-Q�b�O_Q�u�i>]n��#�V���P��)nX0v�"a��(���Y++�Ƒ3Q��

��G'���jz��-��ޭ@��ѹ�0\�f�ZY��oO�_�N��M�:ٞM��ˍ/FV���{����1��{�M�w x���,�X
�[�����;�UB�ɥq��:	��s��� �aX������-l�Y��V��dgnO��Ŕ�:U[� A�� <uG�=A���[T��1���>$�q����Ml�Y��9n}�S�6�3�ŭ��-�-@A� )�R��v�i
i�a�hs�*�X:00LFz��\>���0��^f�o����	Hg^�cSm�I�M���k�L�
�Ө�a[��X)��̿CT���5�����`UK�{HE��ij�t�R>ޛoҾ���$_�8�=_��}����6�m�<a�2ײ��M4��k��ULj��,��E2��Q� +��pE^���c;�k�C���V����p98��!�k��'��ݑ�����
�����J�~=��d���ݥx��6������{�JtU�~T?�7?�����s2�|3�8ιGY�<xuT�ZȬ���\�{aff>�rO^�m��-��T�12�x{�����67wW/⪤�[ ���WM��N��)>T�2\��,�L�}��:Fgx1eÔ�sM��]g�vuhڰ+��� ����K��\�Ww�	��Y�?4� ��p1��a�ڸ�w�Q]~��W��j���d;2�����ƛ�6^0��*�/����0�Q_�w؜T��p��WZ�F0'��2��Z�����
�B�hA!w �� ^�� H�-V�~�ad�ٔ�W�
��7��1W�5���t�����:�.q��~M8����j�f2��65��R���Jܬ�4/l۹-?�0
F�R7_�V��2��z�[�[��1�7IǇv�V!)�T��O���G%n�ѐ@5�e�A}�^0*�O��"�6^5���9�CqE�6*/Уlh��m�u�r�s�	�"E�ٟJJ�*G_�ADK6QS��<�%��l���\|�y����[>�c��{%[é=�e�Nu��R��,���F/�� ��V�h,��CB��H�`��kPW��UK%k�q۩���(�MVЛ;dG�Vx�9@����R���S����\�h��W�V��m�$r��s�BHn.���k�j�w����� �^��>B��2t |����cW͔X�����V�٥Z���#raj��>�3j�6��{�t`{~�u��GJ!&U��v��̀T�)��R�����߼u��o�%9k�J�*z������G��4��eS��P����([.���=̬�-<�e�s�<l�
�3J���I���W6��٭p(�-l�=i�p;�
�٪Q�e>_w�&��|g0���A����?R����OЄtET`��k�%��#6��+����%���Я4X�ǽ$~�������[� ܎�]g����h&%�R{poȰ��*�F�~m����#q<��w�;%���|��/vF�!�˓�����}�����9Wi��b�:�HY� U��[8�憴ֶ��r�Tz�]9����l,/�\�c�[�s V��0���,�� іʤ��������`�*y�O����U~۟#�d���ʺ�+{:+R��(JEM|�v"KapӅ/;U�2Uْ!����E4�)��B��Z|k�+o�_�5��P-�����N�F�Dq�x?��hZ?OƠN;�_u'º��a�)J�5`�і�v	�}Q�}��x������-I�0�Sc6��пj	���5��<�9���
��q�q,�����G���H���r��~��Z?Ƌ��n���q��g*O�n%>_⾦�d(�cJ��>�	o<(B
��v5'�-�˗r�z
���j�@�trBW����'�^-�α�e&N���#��Ǌ�*��Ҍ���L�*�[�d:K3v����c��� t����:�`{�8�G��w�`B��0 W���1��}����-o\]����Fu�N���yy���q����68,��)f�C;��Nnp��`��@O��I1�@(.���6���!�4#�A��n��N��0RW#�[&ӯ��{#hoG��n�q��[�(����ι��mO�S��.��lɳ�������F^ �G��{T;��`���0��R��]��8���\q"�.����a2��uw<P�d�O�H٪)4њe&?�EA��*1;�Y���'�l妿 �|�^H�*��	.33�*F�bwf.H�F��k��m�Oz���s{7�8����s_f؀�V�����[�d ���EU6�}kH���=Ie�����3�E�I%v 7�ÖXP�o Y���,�Ǵ}3L��a���(�q��\�C�C���n��
��n(��?����0��+�WwL�meRF��&���czь>��H�x�/�
�<^�����|S���"k+a��ϋ1bA�R�b�s����Z���<���h�냘����k��+E�
n� ��:�~�$��NL�)���	��V�	�o����
��n�W�t�Q빢-��-��ǫ:-n��
�bމ�	�d���rU���7��,��ZѬջ/h��_�c"e�����&?y�6/pÒ�>V���O[������A7����k�:�HgN��=�rj�}������}��JY�OT��h�Fd4�a��jt�m���N��թ��&�s����f��yfg��1*�߂{��x�O�ϓe�����<��ȳ���[����3�:����R_7�,�w	����ͫ�w+��4��+��	C}��*QD�Ot*w�
b��׍�L?�*�k��e��.H�!��e&U�߄0و@N�D�������,����	�n	�ʲ���zQ37����<��cKuI~{����T�s� �����?�;!lpT��v,����&�*#�)��	��h�����[u&j~	��/T'y;�,-�u0k���u����3$&������0�|��懆2}�Ƅ�h�%^�9dΠ�30�FB��9�޼�wI�×n ����9���okf����gḾA���m����zC�"V�YV����IJ+�3#��z`/e=x��lV]��K^�b��pX:|<���m��|�H9 �T���q[~[D�.�׾�rj$o��~:��vJ���9���	ږ
P�������,�@�>��
�0o��(�w�$O���ړ���.�V&[�ۅN{�m�nn�}��U�:����f}�Aml���/o ��e��>Nq��|�n*��1�c0��sXڻ`��ᄗ�Ts�G�]���fV[Hʞ$Ơc��*�$+���J����K��ַۤ�Ud �6�B8��#���(|��5�(8�܂�^��|g��}���"}��iW47�V��l�tF�I"�0����R��F|�0��ň߶� ����sP�'���m  eǅ{)6Ȁ�sh-�_}'1!��N�K�U��f�n��t���|/��mZ��*4��h��3o<bY!�ΘPb����e���Ĵ�p?#;ɪ��
�n�϶[�����};���wu;�f��
~[�	V�~a��x��'ɳF�Tg8���\���ZQB0��m	d���r�H��R}�Trm�;u�$��vҢM�W��v�7�>����4���\�F���!�𙞵^�nn
�K������ ���Qp�c3,�zvi[�u�(��|/���yEp�6���z��mj���ͅV��۸�{���*ǣLٳm�TX��?��¼�u��|>��1;6�k������>&�ro�{R]��'�a�����K��+�#ׂ��{�X0C���C~-��6=�M����|�.s0�Jz��|����וQ��E�/�g��n�=��4��j��9�lϩ�B�_����x�8����+�m�3�CO�S��:y5˲��팓��L�`���F���v�j��V����ͼ��؋�{D�P��b�s�����7w�`�|xs�q�����͘��x�'�(�@���PU�a��9�rz_ꋧ�y�������@{q�<p��~|�^��O�r۲|?) |{	�����B�汗<%�����ڧ:n�Z�˖��mdyୢ�S���P����JQ�"=r�9̔�e�ʵ���E�'ϛ︹} �uB�D�����y\�y��9M�y���Y��(�.���S��U7�m"s�sH�G��W��z��w��nz,�G��r��X!з���'�Sֽ��>5_1�IJJ(��汽9!ݢ;�D�V��!���^���Or`�����ɳ*�<��ބ�-� ����h�\a."}���k2y�l��9�N�X�+��M��-Pfj�(��{�-I�T�>Ƅ��;��n1�H�.h��+��91rm��Ϋ���09!�Es��.�>�>�u@O��*��X|E���:�r����f$�R7�7ef����/��C�|���JE�yԪ�Nxɠ�ثL΢}��x��`l�m��DDp�N��}Q��g�P�U?~|�^@��&�!�F���/*�s\�v���ŏem+���J?�Tn�	6�R�g,���{�R�Zǫ���┹B r�������D~��9�|E����>�oVVG���v�E��������{웯�]��U���7斝ڒb���v��x@���ҽM���g����?��wiV;��y�����,�+Qhk����w&e�Q�V9uBqN��s>&5����۬��d��5Q9:�ܸ�Qg�As�F�Z}�ng{�*�H��ʫE�߲�Zɽ��c���[�Y�붨*����i6{\��~1mz@�z�����D��[����l��Z��ff��{z��S#s^E2�"+�'��r'�eC�lW�=����F]p�O�oI���7���F�0Î5���;�!�
~'�?���Ȭ1������"�ߔT����Df���߉Ŗ��B�"^\}C&(t�}z\���X%��fS5vR�l��ԯFѯ�N�k�tWY؞��<c�E�g��}ⷊ~Iۍ����[2K�eK�$�\_p�c�c�tW�U�9���ք!�9r�́(U�ѝ��u�=����{��ӻwY�ۜLg~�n�d�šw���$�{|�
�4�9c���Q���&��{՞��gw�Q!�eC���/r*�u��:�l�qO������PQ��Oٞ�Q?k"��OJ�ʷ�k��=f*na�Jݻ�9i;���˛j����cc�n?$�k�EN3�e.�BOq&mw��VV=E#�$��Lw�EWϸ[��g��?

��?�#/[��H�5n�p��^�"���^Vu>)�����M�S��s3q(�_a���HA�ipm��䚴� Gi?t߫���#n���|˖/�DU�����+�v���������w
{�`^��'�V�G
�'|5�l~7�Mt\;����U@hzZ�u�H�đ߰�Q�ѕӤK�X����2�d����"q��C�8�@�9Y������m�p�<��r��Ft����솅�M2z�7Ɓ�L�ЅQ�\TQ`��y�]=�>���>�9V���?����L؇�����/��J����Q��Ǩ̗W)�>Ԥ.�椏g���93*��mX����+Q����������I��q�6���uƁ�C'w�`cz�!u�wM��	���n� ����������x��Oֻ�w��=�nT�=���J��k�L�Ī�!�������}Շ�l�8�~�°�).���氮6/���t��w��5��/����޸��������Ӣ7�Q_S&K5���*b�����ǋǼ̵Y�;�����9Ud��`V܉�[�j��g�c�.��
.[��[�sOڮ:e8�q"[���]�nh�YuU�O��6�p�|:�؃{�v���jp���_�Փ��*�sD�ic�9�^�P;���s?u�	�Ug��{��E����l��w��V��8��ɾIvp�F#�������ۭ�߭�K�����ɠ���[�:mt��_��*��GKv.c߳}
��nc�bO�t�S��%��粸/7'����E�rϏ�|�}�(2P�;�H߃��^�����B}E��ĶV�r��,<�Ǌ!�|Ƶȴ�O��\3Ӝ*����:�I��4�h;gU�ŨE��;�� 
�|:,��C7�<˝8�sW��K�Wd��=�gc�[��$�Z����o��!� ��
��>�'	����-�F����la��������e^Ըܖ�wV=�f�9���C1B����Y\"ԃ�c���2s.��Ws���E�c�[���H�4����j�0�bOѸ��Ζ��d��	����݄�����@�2�~"�}|��TF6���q����λ�Xj�=%���6B쥗�_��Ģ�kd�&�쩑7o*R���;*��ۚ �=N�1)ǝƽK�(�[=}����׆[������q3^E�,��t�\$��D녞���q����{�[� Y�K6� ��$���	I�d�~�뮜��|�+��2�ISa9t���z��7��v�/'�C���x����p!,�7�����~� �V��%�iaI�"ZL��E�9��W�}�>"򚥀���� ��ñ���6*@�����r�G�￳)Gz�{N�٩\�|o��hU���X��5Yrw:*jU�z!��������"�`�8
#y��6����bW�t�T�c�AD��B�
�=�ŃP�.+��WB/�5��E�l�	��`余����W���Sz��_�j&�+@!Hר�nV���J\�՟O��m�X�0Y8�#i��闷c��T��;�ʗZ_ܚ�e�I����M�zY�P��:o�FWP�t1�޽�����EN	�c�����}������>ϴ�N5�W������Ɨ}cG���sYE��sÔ֜ցa���������F�6�1�Ћ���M���ĂA�_ڥh���5��|���΂�S�yd_&H��̛
d�;�$�H;*j��.�7?������='�[��<D�qB6t���o�Ԁ�u]��k؍��ջ� �|�y0�����1�J��8�P�h鶯l��R�?v���O�8]U���$t�$��%N9�\���G�B�ޚ���h�8�W�Üj�6�Ѣ�df�J��Α�����}�P��}O��5�Q5S�'N�K6�<q�v8 ECJ("]�����K�n2V(H
�dU�	��m��,}(�Xc;5�XB�ɴ��Q}�� K�T�{���k���${�$~��];-���JF��tN���=���Jv�M�v�HGt�(�"���ⷛX�֮O��ԉ�{}"ۺv��	:��N���� h��%0i�6y��]M��+P�S�k�A�Y����͋��ix��jzݽ����l��k��A��9[`�Y��Ej�^������GԬ3�h�����CZǈY#�nbD�3���)�X�-Q��$0ʾ�}R��e�WUQ���5v���;�'��q�|~�͎�ћ̷'����P!0oZ�;1Y�����<T(�������f���K!�ֻ��WKW_�qVI�S{c˧m���SO稘�pxm�ޗH���s������->�����(���*l�l�����qpQnk"u�(���X�x]_���g�?�sQu1�)bս����Z������q2��g��.G���{q8cb�;9�$��I]9�E�7~��b�^�l�[���~����e��;���Q���<�5{�W��]���Ѝ�Y��lv�x�<���]zW��XFW_�M��NG[R>[@@�D^��at�
�;u��1+�� �;�����%�o����35̱��C����Ɖ�w
�Y׍
AF@��Y Y��Yx�2:f��Pa�֖q5<,,��իJ-��333����9������!s��U�g��N���Fl���4�q���ۗf���?�݆�I�t�KI
	\��R�u�(�%K.�tnl������<�7?+��?����o�+o��blKђ�Q�ڱ�B�3���7]]�'�L����
M�k�"<���,8��̢�?�|�)�<p��WU��U9�3�3��^C��3����HD!�M�ЌC������n�g[s��]��s�r����@]���G��*nvvV���EA�����N�S<�K�;�bܱ�������&�Y�DTЙ�R2	WS>n�E�������7ɸS�=��&R�SpLZ�ɧR0��m��ݻ��fV��<���i��o!��0��8k�Z���[��.����2�bH��i��ǰ9]��E�'����H����WZ�E���"ݖ>8������~���`wm�������]���=��?�p��%{��	0�⥿%g�=&�z��ܞ���#F,]m4�#�!�r�=�">m�cIW˂ǯ�vF(yix�HR�ZJA�w�u;�U��	�C�/0������J�:����O���󕬮,ag�����@�;+��^���"��\�!�r���n�Ȧ�w�ulQi��9�o�Et�vj�e`�S~��W�g�:�,A�*:�7�L��:��6F�*ˌH��6��K/NL��Y8_�d�z/x�mH�_���D�<����+'��ͭ�~I	���OO~"�=�$�����|l�Y<Jކ�˫�P�<���d�&-^��f�F"�G���2Ŷ�
��@zJ�#ۘ�1��0�e����nd��##��c�M_[�A�L�m`���m��X:��I1R���1R�фϕ��Cc]�9��	�"�����^<*��tzXos���n6b���u���8V����ٜN�liXny4�b��KAGX��b$��IPrg2P�r�G��fW!P  �'k�Sp�S��\��̚G�_�0^$�%��[���(��,+ĕR������i��ٽ�0�(Ai �7lM��:2��*n����ב��KWG�:W32JEWz�VL�Lɿ$�!M�C#��A�ya��>��b���߷�N;+")e�(���A<ϳ������� �}V�K��C�ԇ �HDt���B1�ƢH&C��?���2����Q�Q��Ӝ?F�R����]l9;u�����}5�Bф�&�+�D�W�!"a'g��}�n����ӭ|ǳ$e��m�>�ܞ8�N`����*���M�i>��]�!��R	��I��{9��Z�aw�ѫ��DE1SH�y	�;\:�L��������W�T?�A]jxY��֜�p*]�F�@�mc��ʏ�2Z��3�}��X�X
T;��M���!�6�U��A����v�;��+�5��g��o����4��T���y*˴E�?a��-�c@�l���|,c���i�}_��{�u�=��� �<��+MX�4�m��<��R�bT3��F�F���]�g�����Y�J�X$Q<��Wx]�;�n԰U�^�P�(�+g}�sN���X��:'')^��7999� +�U=�|D
�E�p1��>�����޵NB�����(0�C��ѿ���	��H[�'&���3z������X	:MH�k�J��$��?�؏�A��J�{s�"����
Y����.�ve7Y`E���%��J5�0Q����s;���'n�?�X]RIJ�j�@��EN����<�L��[V��=q��y7:�!8L]y��T��db@/�H�?v�9���Q�eR�::hU�n�ؚ7�:6T��������w��|����Y��q`ʫ�A�"}J�:H��1
���l
xD�Z�������y���;s%�eMX�G� $	Q�?�ev��#`hE���,p�L3_{uErF"0�yhJ�%��
���0r`����I��~��=��!�
M1j	eR1�h:��]��T�a+��2�� ISqF�>�$k�84�a�$��߉43u��"��L�R��un��e�l��'d�Δ��,�9C��^3����~I[}ϸ���~�e���I�H��o�Z)Qr�v���	-A�/,�8O��k��h���z
�⾱c����k����{xʱH4���t�|c����h�)����ѸMQwstZ�A���	���r��R���zZ�U�����w��!�������
+�4��qm��U�M��\e-P"���̔���p��濰�袥��)
��t\I�9��R��=q��4Y��k����x��,�02�a�g_қ�k�� v�Xq�0f-n��ż�y3�5�Q�t���UV�1�?gB00�ŗ��3��cLmP����<�>L[	ɞr�U�,��"�$~oI�3�뾘Zr�:J�3�8� f�P�M_7DY�:�e��!f|G�WTu�X9f莣2	���M���M&rؔ��[v|�>^0�0p7�a������&fmHt����M�j������>ioե��f�5��Ε�Wx�� L6��t���}3�a��-P���
l�s�}4�i�՘���9�K֖�mOY0���w3@�6t`�V�ɳE���Y����������粲�O�<r�@]���E��S:�Q�]9n�!����q�P]x������ꘐ�O��Q�(�(��ȯ �0:��с��u�D����B��d����H#���,�'-��%�n���}n�Yĕ�뭉��ڭ�L鞻_'+��ZP�N�����ҁ��9���	h����;t5���q;b�f��q����s]�h�٪3���y�M4��u@������-o��K� �q��$��ǢsR�
A�})N�_!�t<��f�"�$�i3]�����Qi�#��b����]p]�$Z5���+�FR��X5�4�n/e�+̰}.��1�-H� �����;J]!i��B~��z�t3;)+��I��^�Y�\��謩��w�.l�xY,Cס�t�3�	�t�L�g*8�Bn&~��H�t*O�حv�-�;	m�|y�|鐽,�n
Ջ����T�[������R�^�M����C9�.*���6��&̔(�ZM5� A�yd�-AG��6c(�&� � m�B��T*��S����I�o7UԱ�5�� �̺��ؽ/���L)tZ�/�W�f@���=L�Q{�����w�@�K����,饪� �-Z�'p]�,ޏ�����k�:e���d>����?�:��"�H4M��y��GN�Űr
MM�w����S}���++̛;!p��)���&?�4�Hd<��uӤ�V�zd�Ec=���A[
�Jݸ�����5K��:�2��6�<ۜ�h�5�iN�U�n��]+����:~�;�V�$����so��\��N�Db^?������l<�0�����xFҀ��`�B8��%��d#��2���8V��w1��|�c7:�
�����T�v���C�A��	CfV�%�� .|�D�p$�jI%e>!��8쨛�B�p�D'R<��W<�+.m�(Ʊ��Pq�C�t�������	Ȟ��ʝX����B���?A#��WCg^+�	_g��N���-[{���I&BP��W��:��"�Xʹ;���	��Lg����`%aO5�%}V����EMt<�����Մ�o >u�Yi��Y��]�~!�m�[�/�VTv@�+���s�x3��G=��~�]UC反a��F� �' .��JT����W�wT[*��K�tlq���g\`qy6��u���m ������NZ�j����[��\A!	��d����
<�݃���UcU.xbhS�g�!���9/Id=ڪ��GV4�2Ps�R�?Vf��r�h���*=$o%U������ �������L(�jޑGKw�Ң0MPnsj��w�B�_�<nz�;�n��tǩ�R����xK�	�)Uu��DS?��~�H�۸@�s@	�s,6�eR�w��"~	&G�ѫ���?���:�&[�����_����@�������Re���bȗC��,��a�Juik5�����{�/}R���=1�&G��>ٸ�aJ�oe�M y4OnA;��=�q~oe���7��2v0&S;���H]k� ٕUŴ����<�'M "��o0��N����s��H�����<f�JU4݉
>��u�����,��^3 OF�tO� �@-���J篞A2�-[�MI�J"���$w�MGE�G��0��jVYVV��Ɣ�@ϡ�T`LW^��0�[�'@dd����� �E�c؝P�o�Rd{�Z7>�-�`đ��E�))R���+�����M�b�B)��ɸ�Q���|�d�FD <��-ѣC?!��+.&m+�%n{�쑵*8�9EOB���)V�B���"Tu*놏�ϐ ~:[25\���K�OԒ�	��8��"����Ͳ,��N�YJ| � ��,�V��DV�w|��h�ʮ�2��BM��7�)S6T���\yoγ�p��$s�|E�pO*[�ܞ�����}U m>���s꿉���=s���{i~��G�@�|E�;�^m��qq����#��4f�[90%��h�E�S��bn��ך'��g��*Ͱ�����������w�g�~�y��fʂ��;%ކ:���5s��[t�T�f�4����<E_�\�/n�w���3��1F�+5�4�� ��&�,_]�.�/3Q+^���N�휀�+�ɇ�.��!
f�p��W}O@�H\1�_e�;�o��mi'�Y<��AeL�.��8۝��8KW�A5~
`���l����:h��}�:�c-Ge�t^��4���e�GHj8]i��L��N��=7$���4�Gˬ�+#�+�`
tu�D��?��h-y�BZ�a�ћ��5�RQ�	硚�?��hj)��E�$Q��1^�8��b���Z��;\-}�<vfey�Ң�á�>A���{��AgZ��,0���-��)ALsJ5�c�o�ѭ�����&A�[lc3������f�,�)�ǎ8R������Z'�y��뱨�Ȼ�5pX��X��%�p�U/m;�󀦂႙L.@B"�R�z�s<
�ga�]'�B-�&{̈�N��G&�h�j��X���ԥ·�v<e�ֆ���b�d��)��pr%1�b=;˘O�r�R�u����]i�T���EE��&���¢�:�~���������|��B��I�D���nI�����I~���~��j䐴Ïz�ݟ�^b}�"��=2�e�� ZRF��"��W�1c9$�س��qzV;	�u�vj��*�@�.8W�
�;:�o��	�`���N�H.�5�5Y���J �233O��S��GGG+�Y��)w����拈���(���$O˖Y/(��g|B�鷷���_r2 ��7:�=5Կ@�//�4W��T�N&�XT�
<��ZL���?>ca`�8}�PP����&��:��A}Sg�tE�@w9	JՑ-C-i�b��I]T�?���!�/�Z�)�M�rz�"���	Cú<S)vJ(�sO����FjG���+Z�V��m�Giq�s1*��1\�X]̘�lj�:����o�Y��N�U�� ;�Γ��\җ����4�鿵�ik���Z'K���F}F� a\$w�� �ڙe���������Լ���pt`�6ooV��-8k�5�\5�/����?��_�C�T��R#��"#����+���|FP`X"$¢�I��oO��t�h4�z�҄5�{��_��N��gq6�j��nvR�h� �ϳ,d�9��ϼ��vSR>�����;޵�A��*�S6$mEp�Ei���wQ_Z�$��]�I ���;�q<SsN
��<�"TE������f� ��.ڳ�Z٦�t�"qP��_�o�hr������!NnJ�DwY���d���ǐ)ޥ���@&�٨�ɯ/��y�UBҐl�܏��~5aW�E|/������5�V5���h���V��O�t��VV����w����D%T�I ��Y��3WR$:l���k(�
g��:_U��,g ��{V�m�U2���iа�����۵1]�x3���y�?:[]xeoP`��;w�fG.�n��B��L�#yh��`�s�bH��S�o�H�ΙDgY)�Yy�U�l;?����T/1�r�oZ_���������C%0������^��i�-��^ӿ~5�O y�vk����w���Bժ1j�I���#�"Q�}��U��Z3U�V��0r�S����/�I����'�>"����)Ԯ	�r����/D�J���)���1 y�у�54h��7�C��m�3�B�A���k�����V�={��{=��S�u
)���
��J�E�y����eן��fs�c��3��)G��"M��T�Z��"!���q������&�	m�f���X�����S�ƴ �j7���e�`��8����������
X�8��-Ʋ�b�|1�9L~���˧m0gSD%��Mݴ�E��+s�+ݙ8�E˝y��)����H�H�Q		����`;[�m�R��u(��0��a��[���fflg'���͉VSݟ�wCv�r�㲚��G�$��T/\w
�^Z�jrEM��v&m�����t�-6��9Lw�Ug��c��G����0??a�;cu�����~M�U�3��?x��%��
�xx�ă=1�}��GQ�vamڃk$���x�PL�Nc���ft.d���:���u�<��*���(����dK�g;��&�ͧ��#�_)j��}JQ��J}��@1��H^�.��V�݋��8�t��T���l'�����p�3�4�:�t�����Zaf����3?��A�(���d������+�;ǿ�/����ĘF�!U[���j��@�;e}%�{�'�)R��W�O�M�?e,H����wNm�����_���O��㓋<�{Y�{�;;Z�G��-�M<5�m�3#w���v-8���{�RUڹt�R�D�[�!,	��a�O���&��x
d���� ��Ss���a�i�y�6��:�K�C�n �}v��mu���ں-~N��j�D��mn���L�O�7����h&v#,��M��c���QDZ���j�a� gr�{i��5�51��� �S!�fQ�<���u����0��jK�@�xos����O�Ш�<���_��d�t�����-�P�h�&��ƂΧ�$]�=}�y�P�����u*�P�Śx�Ζ��&�~|���8w����[gg��g\	C]	��L�$���y�*�Ko_ZZrpv~8�]7蹏���+Ղe5*<vk��]s�@r��Į�G�P��'D=b��Z��u):8ςX�hg����bhqixxx�t�}n�C��!9>��\�|��-�;���a;�G��WWN�ċ1����=�`���q�����?az��	~h��+�;�F��ɈwM~��q�����%�O���(+fq't[Q�@��t�����G.�U=�B��<�������T�����B(���>��j9V��W��� �&�o�ɱI,��G�O�� R|�Uǖ��[s}%�,\����Ӝj�n��* v}l�����t|40�	��Fɫ�����d�p7j��3U��0��+UYs�y����"jVvr�	�̰�|-w�h�ͱ��Z�.��l�ƀʚ]�����)��EB�q��Q?�!,��+n�:�����:����goBo%�ե��xJl�����m�6 ��Ƕ<�e3���λ�Y��^�����h�N`��D�;�`��hC�
�����8{��U��hv�;�i߃E<�N}_'&@Ş�R:,����gx�+Աy0U����L����+)�|�Ty?(\9R^���P��W).���h�p�˞�`���~���U�B��Q@���}v=i�9^X��U����	�5Q�6x bM�?�5Aݸ�ѝA]�e� �mv�X+�8t�{{v*E|g���E�G�`��㊄��d4۔w��:ZK�5�{����۷�M%���V�*Xa����	زo.�c�[�c�@]R��TJ/�,��&JcV�~�
iڻi쁅C�i�z
�2�h>rX&��譞AQ�R�R&�@��LWvj�P�(�}Ud%�� Ժ����VM�q���~�*�@�gU����P<�e-Xek��
OvC� u�J���;�6r-��Ȇ�%񆋶�g�e��_lb[������ݵtݽsnm�����L��i#�'v�Oa��YFA��Lsҧ!���(B�t�ߡv�4�z��Ӱ�ɷ�֎���l�̺��#D񗘵�Av�@V륻
�A-[���Q?D��?2�U�	�푤m�z�'��߮HǠJ��?�X����L���ae��ARQ+Q��VMX������N#'�jf`�ß���(ts��)�mA�%���<J�N4��EH3��j�����$x!u��L������9�wvl�IC�K�	%ܢ_{V� ,Qe�<��hK�n��B�'(=�T�F4�u�Q�`��d�r�J�a���b4����8�7��%t��_�%�������k^3Uz.nn~bO���dsfs�>��YaO픆�ϼ�)��%�uSU�,��=�Egm���l�G-x�jN8�uu5��2b,���}d
����PC-�L�b�~;�6->�v�~�:�S�|_���ͧ���>&��"��ڳ�"���5��R`��Ҳ� ����ѲP�l��
��B�`���6��s�5���T��f��veG�s>�6�<�O��7�*�?r��J�u� �O���1�}J���He;V��6�؎��Nͷ&>�>�Ȑ�4,��Cђ�j�/���
]aC�;�*�#LU�Uq��i)3�3����b��V]�̛�>F��#�k�Q�m��"S,�!Za������ݘ���iJ$5�."����.]�	uT
�zҼ����V*?F�T���}5HW�䧸��K�Q���/"R�v�� �s�o˷�w�mh�2�����_:S�s?��!�Ó[����j�UȚ!*�@u7!��9m��K��<7�^�9h��p�g��/��M�|AUJ�|�і!�y7ZXD]��%z��X]�0zoe'�����ԅ�R8���}Nb; ^��Ї=�������{��E��_0}�H��v��D�Xfl~��^����Y�^j�H��G� ٭��z<��6׷ -?��p\^y�&
�l���[�\��Z'��H�B��{V4Q�Ja��ޠ5(��'%������	�}��Sk��jṁ��B�O�H����@]ӂ�?�k���Eo*�3m�$�dnQ��žh�R�ΒR���2�Ͽ"搐\#D�HD2�"����9o!"����������B
-��b+V�������2�6d���m���݅��h��J�,�P�`\I�ࡇֳ��2e��6��Ҝ�\[����`��Ls>�,Ȧ��º�%�M��EQ^�]y�Z�,#�����7ڒr��6�lE��O!�Ei��7�.���{�xڈ�X��yvb�T疟T@���k�o��0H��p�KP�_�SQؖ�E+p�Vlg�-�)H�p��M
��Mjy�lD�;w<1���;!��g�$���|�J"]�s�3 �1D�����Ƽ��|%NS�S�i[�A��� Z���C��U����v�erEE�\������F�zM�.]��1b������,L��Sc�+�W ��JM� 0�����Awhz?u𜧲�we���g/U���I�U<��7���0��(���E ��N#�����?�;����F˟h :��zʨ��C��|�C8h�vC�R��9�]@���_FG/��X��Lwi�£��pR�n�@���58���� �`v���Ⳍ;�	Ɠ
	@�>�jU����'��࿙����I�1��Ko���Q�ku���L���~� ;>���i[l
�e�襕������%/h/�d��	�8D-�e�g�^Gu�˖�e�<X$,pq�@C2%��~O�1�H��EyT��	ˣ�q���ӑ���]:U.5�mS���_�)l����,u_�zh�y�rC��t�kC�w%�_d�	�Qf5A"e�Di99�쩛�Đg�_�'�f ��7���࢚����* ���3 IK�(bOc�$���o�iJ� �J���u5�.g��}���n�zɊ��`*���B0j�w8k�{�����b��Fi��k���wT� 7z�d�Lź�u"I�����).*i�{�i_K�;V~�;��i��ܛ�HS�⻨5~�nn�F�NJ�"��}SC#1�������Qv��/Z\`x���ɢŅ�ɵ�!��J�8��X�MZ�N �^j�C���-O����M(W����{Xq�!�~���JR�M�������k=P��rf/^OZ���8&=CC`��{l�� N��_�ߞ�E�q���[�����kbl�lBw �����V�CϏJ���@.�h6U�DVQ�Z�	n8�{�o��
�ɴ�dF;�4�.����;Ë6O��]�w����*��|2)�=5~��H�m��z}��L Y���3��h����>	�
3ป[��kvْ`���g���A��l����,�XH�h��{Θ�P�ړzհjn<��6�.Ȣ�����T�@o��.]&�EkM8���&'y�sN®�_��G�I�'�a���m0F�����!s�3�;����gZQ��Q{'�1�4�8*6:���3o$�%�>|��`�2�{�e���K.7]�O��k4�l����w�ڶ�eȔ$)��E$d���d*��1eNې1"c��Gf�)�$��B�6djocƄd&���{��{���pt���u��x�����3��f�
nx��������<v��kF�3[RC���Fw���d|��R�+�ӣh���6-;�@�����u�C�����{��*Q�<�T�3l��c.r��_X�ŞJç��w�aAn}���zZ�vmv.��7�:�g_�Gێ��c���H� c���6e�m�R��w���Vs��?�<�܌�%:Ț77~�f,`�r��Lw�,N�5mH*��475�{je������9�/����3!\R��sm���ɚ��<�}���N�x+��M�7��/�^�̴�[��"D,T+ƦO!H�}ࡠ��mL��H�@�W�>=��	�Nǥ�c��.�*�R�)@��������4���8��/��E�3�T4�J%T���d���P�g��ҽg�"�XȐsK'kD9`��ۈ��~��疸)��q����K�g9�zE��e�M��0;�9d�i��X��B���qS9<�s���=4%WiM���Rŀ��wM����m�:p��B���6���pX���Gc��='�#�iYũ2�+�^�QD��|*̈�9�ʊ�h�|/KI$K�܈���1����;ٌ���%C��#�� �N|˴O�K�-r�<�Ǩ�WmT����Z�u�ûj�g����ᨧ�sdu"HS�n����`�PV�tXdQk�i&g9����+���dȭ�G�:oS��y ٛ���bc��w7�g�iP�A	`��G�ٮ��!�,�dMO`��%�!�A(�Qg�T��tg���S5��w���4���1�[�ʤ�=%�b���@��}��Rb��g �c��˓��^;4���aU��̔L��RS��j�lo=)Ụ��&��Ɂ@4pg�hp���Ld�h�����h���S�eV�����2F�#���RV)�n�r3���ve�5�HEԾ�#�ݳ^��[��ҴҌ
i
U���gL\v"�w�H��kV��� ���#�9Tt��	�Y�X��]"�)=-���P��">i�;�������H��U}Z��n��w=��c�Ýrw�3*�1mr��ie���靱�eGN{�j|it��9j��j��~�r�`d��Ś�P�'��<��Ŷ�-��z�ִֻ�;;�Z��؊�i��}\A3s( ���ҋ���V���'��ER=���r�&��QI[�ee�pG���C;f9S���H|7�R�0����U�d�x�ay��Ԗ/�Imw�ܓ�0��!�!A�����(o��Y��;��}�PMfI���.%��0+��\0��v��'/��(�[`)֬�C�~j��n��4�<�{Z&��rCC�ÎB��!��,j�O��IR�;A��h}3)����7��P'�\	f/���+�@>��ߒ5別β���&2p��4%�)���BQ��?fx���ϤG��L9��u2�w|�����Uk����PS��~rh9Aj�p7vN��[28m��)����ӕ��ٯ�
�����,|80V��;Ggjc�ф��|^{0KL4���Y5J m�ڀ}����G�C�&Tܤz��xKX"�h��;r�NfZ�5��a��e�s4�5jK�A�3�Ks��Yb�9gj�><�Ƒ��M�I]��Ȫ1�� 2��{}�Nb��>577�.Uj#�܉����[�I���/� �f��`Q�9�և�M�,]cX�%$�tb���'��V�3@2���]h�,O��N�����;zk[d�eT��T������`P��<y@g.�t�����[�߻�@KC��G��3r�)�1���=t!	���ڡY?�e�c�G ���v�f��Ɍ�(��l��B����ܔ��!S��˓���HYp�8�oOk%z�+���7&��N��(O�B����K��>�i�5W԰�-����͸�uS��,G�T@�n���4c�p�)��[�r���]�3T�F��� ����q[�ݽ��ژg4qeAN�蘭($�w���B�C�Ю^�dM�� 4���SRݢ ν�ܳD���v��'��ͥ�2�)-�����ߡ��R���$	z>�K��pB�@��=�ҳb�9[8$o5/ ӅW>������j=3�d��v�R�˽��.a?� v5��c`��B�~1�Y4��|J)nA�c�[M6{P3=!s � ��h��]���E��e.�i~�T�{y�TV��PƵ��8�q�-%01@%J��u�aOK��[����=��ۍ��S��*:�H���g��vx"�q����8�VF��1�����БH��bǠ�vO��������~r��5ܕ�>yz�*/��l�t(=rx�|�|�'#_�B� �(`���^�K��jF8�NS#Wg@#;r�J��!�v4K5�'�4*Nº|�[��e�Msu���ݚ��Q�?��y��9�< �Ա���S/�	��E.pz��1`PNMۚ�E�%u777����~��
�"<�Wr��f���%�W55�󋋎
g"6��o���ϵ���Cz�P�3|�u���~�._f��������oS޲��5�����SP��Q.���^-���r:g��rd�3���Qp]�Ӳ��}����Sy=���ǣ5b|}�����L���xiz��*�$�y��{x{�gd}���3��s�3�z�@��ʭ�p�;�1�1�(|�pX�g��ߌ7,04,�TV.5)���yqq{{���`��h�/O�om�ib'�I��c�q�Ե��ƽvp�CEa������FU9�sY8c8�8�����)��ײ�.W�����}��K�__Y9��L/�vA�(-ZY�h*�`��,t4�A������!%5U~��s���@��2�Q}W�+�+Ⱥ�Q��yO���L_7�q I�ȸ�:���n���7#ߧ�D/?ۧ����w��57��V���A�H�Ǐ�O��*ϖ�?���1�S��T��*���`@�;�D���i�<rP��ɝm��bc�y���>�k��e�bc�b��S��iu/,�HIKW����P��myϮgDb|��}�'�#:�D�c��Y�����2������(�c������4$���Y/]O3�-�_\|����p�^x���kA�>�����oA�v�����ّ~I
?��)�p�6u���ʔ��5��K�*w�W�:S��V�֖�aX��>����S�zU$�;>�-4ڱ�[�)/8s����U�ѝ���j�L�8�-Sog:J�*����U_����s>k�l�*����Q}�����R�C��?����\Gk� ���C��{��
�P�{lea�S��j;�����Y�9{-���t���*�v�x��p���W�����\)��>S�������������7"Ѱi�l�j�(�Ž�%�EV:,��kf��Z�%��	�z)�p�����v��f:o/q���(��YdD���K$�A��ҿ���SI)��C�)*e�.b�-^���2���^���0���l�ֱ��a���	�=�sM[�ݱ���=%�҃1-[ڲJ���b��V�}�<���f�X_�t�'\215�:>�bm}*�Cl[ݗL�Õ�?Uh=��ym�]*���&�E�\4��5"/0R
2�}���^�ۙ���7;��C��	�����Sԩ?�a�ܯ6�u��#h^ʍK����&�}���А٣�zj���B��d���N���~��R�c����˓y�,"�}ZB�F��o�5x;��&'g�o��	�J���..)A�OVh\Է�YU%[ar~����5xI�\9=�����;䒺�.��vm�iU��Ndsb�6���֎�+eO��*���O��&i�ǥ��j^;ֹ�I�x7Tb|�Qi��:S���.o߾�1(h�T�\�y�"���.�1��B��jA��|��7���Z-�u#���9��\���^E�(|y������ڌ�����*ٝ���I� ��C���/���&=)�|��y����V��.����ng�۴��#ke�kd�ˆ�<~� ����L���n�d���eG����%����k�**	��V��s�~(��1]`\d��2�I���2(4�,:���j�n�8��ڢܗ�M�<���_�i��gU��KIb���ϵ�g�Un}���cv*�{�U=Gl2���	�f�^�N恔>��L�X[[{˲\����?ۤ/ԹԸ(�Rqp��j�Io����`��6���U�×���?�P����N���ʓϏ�g6����L鱀P���M�z'dS�;���ܗ;aTd�h��{�������1�{R��0c�3�N's��2j*���Ǳ�[e��f���
��?�ea9��4�݆l}:�9aQ]��>���Ae$�\����z�v��jQ���j�;��sײ�gT(�:��I�x9���C+��T��m��]c��9Lvۢ��^�'�ܿv��z>9y���+Y�)�0���fuM�_d��9b�s�Ǐ�5�(WՖx��!��,.��	$V[e;��?m�Z�K���K63�0��+�cHuݵ���� � \�ЊS;�I�{�Zo�i��j|z��Mf�@��G��������_r1���rnSQ�6/
��ҳA}Dk�u�\��
��[_�s��������B��?�WT�oES�VNQ�0�VeF�o�ˑ,"y<4�'G�{*P��ˉ=��Z�Ӵ��9mQ݆�^�~�:yIPxi�Y7��[\��kN�7��+��5���ږz����hi������V���P'����\Y���vy������?ߤWhʖ�{=��,Ѽ��a���^��7����(&���:3l=N�;�)����g���V�5]$�l��Q�Xg����nD%i�|s/�t=����J�ҟ<�}m�0u\6i�Y���2�eW{�����S��L��+� ,���א#I�/Ɇ5���z���joow�J��B��s���3��M��L�?!D6�@S"n�%���	H��!��_�|��y3$�m{�_ӷ*�����B��6t~�#�P�� �����뼇:��	�.:�;�چ�/��uV��ǥ2`�&g�p����٩����=US?��9m���u�a1�L�^镑������S��Jc�>�|�9���+w�"ק��7�d�&�%JB,,,�g�sutO�)�Ca��A|��0�zU*=�>]�!BFv�dSt��1���h7]+57�5(3�����FDFH��޼=8k���U�/������e��M�B�$¸�Ky'vM!��oJ�k
5������@B �J����j����rD�@X��u|y�MC���ݻ�67��������>����ã:y焑`�WglEuu�`4{��Wz.�'�����HK'�pH�L�`�ڊ�jLTN��Y�(�JW��*�n	��EW�G�̓���Y���;B���v-��N��L�֝MSZ,���,�vw�Z���!�J��0xB�D���`�����qvvH�G�G��:�^�K��"��d��nS�
�g݁�tdyK��W ��yIz"�Y`!�q>��wi�_G�Q/zhcV�>Ģ#��� 13o��g�1��B���p2v���rڎ���������oO]�y��S��̞[a/���au�>���P�nK�)c9�6|}}���(�O�:A��O}N�ln���?i/�z��
�ٗ��ݍ�_�����QLXQ�Iβ�@m��l�~�[��idg����0Znr�WL�Ջ��w�\��$Y��?�H>���~R�bT�Jʠ���8v��rv��^CƗ��g,��u}r�ӧ�/��������9��у�㗱�#MT4��KW�5��M�0�l���w�r7��A�uk�L:$=�X>�|�2o��)Yܞzu�1�!@��eD�{�V���	��;��l��Rҙ���k���L��/j�Be����P�Z�<D�ޑ�a��e��%Y֙�nmg�s�Ŋ/��2���C%¦8�� �(�)���=�=L����7o������{N�;}��-=�4��p�a>�@K�v�E!�����9�	yy�Jm�Wm���O6�O7^V����P�C�+��C5A�UyPĠ`�GoQJ��A' �2�#U�,N'�^ݿ_�q�vq	2.P�r1@�-�G�P�G�.�j.�� �<�H���4��o�s\��q��!.hm����P�.%C�'I(�Y
ſ"t;n[�o���xy�ʴD �MG&7��{,U[ՙٟiΚ)�]q����T��
<ktC����P���ZX&�Ge !�����7��x׻��w�}��pC�+�G�����	
\گ�9� �_�v������	�Sk����g�(^\��f��117�2̖A7,d�~8���0OX~�x����)�L�{�*1�L�V�
p��rJt��,-W$�&�pfr��)�B�� �k~5���0\�3��ȷ�f?}�T��w��U�V|���1w����:�02	rU�b��0�'��x��Y��hՖt��_��ӟ�Ȩģ�ݎ;�K���TU3;�0��,5���p~��� �:����}5v2�4/��m�qDT�}j2�8D����^�`�ƛ#S�g��\nI�RF}�����f��b?�s�S:%=f%�̀��Q��]��� �6{w��^A����7����5@�V}�Rp
i�#�N�Cm�R��;�'�9�ݐp�ķҜ����^.�K��!�a�Z溣���C�ftXNs�;tK�f～�eZ+$�\�I�z�Zt-Ҕ{��IW�̖��iɝ��ǘ�?m��e<���\7� ��u��d��~vߕ��m�#��B�X�V������ؼPE��sdBQ�[���s"C�YfWwJ� ���ۮ���.Z��XyD��l�p�ۙn�f��yB�N�Ѓ�.�Rz*��_�����9��O�O[>�:�����N�7^���<+"�&@�R($$t����U�u ޓ~m�9_[e^�O�0ę��ޕ����x��	$�=���q��:����5�|7�3�`"�\�^_}{��{����������}τ4�)h���AS
S���ګy���2C����I���`���m̪uQЛ�@��U�g+�-���s�fjm�?���$����N��)��7a��|g�]���?pTE�7����j�5bA�����z������-����Y�� ��2Fd|��>�(��ܞ�$�+**����٨�<f,��mJڋ?6�%�y-��u
	�(0�������_��4�Ax�qc�E��0����{��MF,��f"�^���c�	iռ\ڟ�D��H
V�����sH ��K�$��a�</��r�y��"v��+�v��	7�8��kq�vj{RA$�?<3��/��.D9�ss��H��n���S�fd��SS��A���7���P̓�#��:>PM|�<Xӌ��(�5��
�?�h����y"S����t�3�s��P����)�$˴��^S����b9!���g���պ�V����w�cv���_�n���ᳮ�x�S;���Q�~��|c���as��}�i��JYph��s�a;6��95�� ���fn{K�:��Y�w'-�s���g�!E�1/zf_
�A���j�@'oUm=��O����<�c��3̓v7�C�Ļ�OQ��s�F�&~0��4�///�4qB�sN��-`�0|>�Ξ��]��?�KW~�����F���\<	�,����!�JJ�3�`}�8����5ת�꟭�Li0��?
*�����i��#����m�QOi]أ/|>W�#�0w#|���?�e$�c�T_�2*~v�ۓ�q~���헴23��j����hj�KJ���,M�Gd��͵�[�*P�p�9��y�s>��F�����
r"I�+�)B��:�|N�� !�Z�_~ZZ�Q�fؑ�:��1�5~ͼ&�Ήq�y�uJJ�ŘD)�:<��0���&��>��R��BIP�D�5U@���NmZݰ���]=�����S2��#I[�t��u?Z��B�?��?�Fޜ�-�F8
0��mPp�:�����>\kɍ��'kj��":�b�3ִ�Z@|�_���^�i����Tk�aQ��J�{������+��H\��dz�:�լ�0J�x��Y�rSq��U�]�ku�����]^��"y�Oh\�h�Eٖ�Ӆ�v����juӡw������9����9���6 �P�v.�ꓫ�*��-�î��Tb�*"?�PS�$���H R�cݾ<���n-��>��'lU��#�`Y���� bEׅ��c7P�*�n��צ����7.�~���>.�·d�*h�EbsH8�q,�Ylu�3ܳ�R�t�8�2�D�
)gΜy\Á�, �ۍҾ�Ʊڽ_=��i��ѣG����q���F�h�C�h�W�}�ֿ�Ekҋu�S�%><;~uV| eܙ�]c��|+���u&��@{`6g��v�#�iY��^����J����֍�;�UBk�Xgr)�/.@�1`����
1Ĵ21|yJZL�/��վ��Pa�گ���S�h~�y��-~y��&4Ayr@ǯ�|�#j��9��N7��Z]�;\��a<��Ni���,��m�7�niQ]��nh Ƕ�M��.�|
B#��tY*�v�N�M�ESx��9�P���Y�Q��Nh�JO,������ɥ3��Ֆ{�P�
�m� �j���O�r�xv�E0���Ar�����ɰ63���.�z�e,�����}lͣ�#�3i��47���S���JTUJWJ��Hu`|��w¡h�X"Յ͛�4�{'L0{�$��6S�?Ri���Rb������8��`t_S�1�鴷Π��)��!���j�v��N��K��Q��u�*@M�!���Hy�-��0�k�6��ʆ�ڜ~ii#�v� v�n�j|Z�ts�Z�ki�T7���Ξ={�e�tm���Ʌ� {��[�u�H}�^~�F�Ӎ�w̮�� LD�\��kE��V�7���;.M�c�+=V'=�/���V�K��L�H���`7�u�̈́1���E�֝~v6�'�dm*L�ے[kN�����IO�%zӘl"��JB8�x�q�Di�}�M!�ØX����:G1z��Pa^�+�D���P,��@��J�����hY|0�lV`AJ��:�, �8��`�6��D0A��)���i�#�(�<��	},��kP�_xL9z���P�^�mrӦ��/+̞��u{
v��w¤b�V4�cHl��|����
��2@�,0�q>�*��Q�c��3G#�2��P������z�/
�y�iظKљ�$��W��e��A6�O�h\M�/�?�j��Ux��i��6�,���>������%"��򘫾.=2a�O1!��nǙ�C�!���yj��Y�;H;2�:]5)>z��I�~�F��2���Y��.��B����_*^�����>�=__��^�:��9������	
%� �9j�xmu��Nb�qѩ��5����P�>�rƶۺ#U}�������2����#�7����S���UL�x�(Gˆۉ�<��lqb�.;䪯��鲋�/ٴ�PK��:��J�
	C+d�QY3κ�J�arNlrgmd��gB�p|Th��$�:s%~7�<�Q��(ȕe������P�K=��>�,�>�q� *�U:��z����	%�%=�ߧW� ӈqXW����ٙ��w��&<�T_�g�^i���ࢋ.�y婕��[ev��IZuQQjX`���^�[k9�ǀ]o��9�Ɏ�Lg�M>X�̀���,1�#�䭪��Q=�*3���ߐ�.��o�ܚ_���� .xs��Y�r!9{"yР��s��:6<3B^+E������c����U���8���B	0���9��.wB�,�h*=���	��Wʒ� sG[�=	c�+�;���S(ꭥ�K� ��WVR�F52��5y�l-�)�p�Ϝ1��;�KA�B*
{4/��d�U�dc�J:L,��fL�`����x�U�.)F�.�åׅ
������_ϥ�DT�[��(�2*�
� ν�|r~��z����PP�RS�,�>l~V��8J8��y�1\u8��6�O���W��*�Ӻ��PG3���JV�*����q; ٱ��%���YXWD�,Q���?d^�m��Sk�YfO� j���!�%0[9c+Be��AQ�[Js�:�z�H򧣛�m?���� 2Z��
�"}PCʙ���駎���
_?s����ƍ2����|��7��U���q��F��֕�b��=:ݝt�v#*J|"�#�[��<<=��Q���:�8$�A+��s"s�g����$��������i��$����.^s�[.�}+�7�������TVk=[H֚Ž*���ˆ��!}Op8���?㸧~	�2�'�q�v��%W7��w?b^޻�.�(�8�����ڣ���ޭ��O`�/9������s�[��;�>����`���&gۍ��mS�{J�H��xzu]I���SσA*u�M����&��~�jnȆ�߉�����@U>P��L;
��yfʏ��[����]$�����(��6�֖�˥!����y�$.���|x)R��܈��U�|kE�����`�Hl$Q4��F�x�y{�pf.�A���l����r�Í���� <Q��q�ڌp'���.��#�)���+�>;UW���/��Nѯj��3 \g���|�۶xka��W��7�ג��W�u����O�`�kK���P��6�/��v	��󋆥_��^-�_:f�3�'g\pC��?%���[ܩ|E^��J��=�B��d�X�o��L;6����J��d��h�{�_9�x�%8�a��Hk���s9�$�g��&����T���B^�]�>x�A'��W<T͋L}��������N�zrI�ř�'%�C����IV��{�n��ad�6'�a�
�b�?�a ��l�[8����5ׅ���˷n���
ΐl�%�1E�ǫ��'g��0���;��i�+�J��+��ש�l �	�������}�s3�G;��[�@N�� '����.��a;���� 䑂��մ�`�b}��:J�[^?�Ւ�q�t�߇a
�`ں1���ǩ��Pn�.ݭ�'�<7�3�HKˮ�<A�4��b	f�9�lO�l���]a>Jl�?c�R��
}���B�u^�E<��v�d�������U3;|�RTTDZH�H���ؕ�믂ј�t�P,�N����ᴁnLk��������.�,����R�w�3���m�cX���Y���GKoc}��:���.*�����F
NP8����� �]#�f�gv\jU�"�Ҧ�nL���\k��Z�����Ȇ�_�8��b@*�E�_�������W 8�CF�Dt�4c��&���lc��o����/�!9�ډ!�'\�&��6�Š�zhmqh����������*�W����^��i�˂�/#�l?w�a~��ՍǐX �d��~��C�Z���u���,΋!Y��O��<�[+?�Qi�r�����X�����{��k6 �w���P��w�R��;��އf�y��Z��7��D��=��w䭝ؒ.c
ݒ	�B#Q6�e�jr/��ɏO�ʤ`��(�ye,yB��2P���]5=�
�ݻ¹�R��z�j�΢�۝י�o6�P�I��Z�s3^��)���hŸ�>k?^���>z�$>�x��F�-_d���W���Oȫ��7Q�j~�������q�zwcϼ��7�M��3Nz&ƞ��ۅ��8TC�k��+߿%��̶µ�ґG����7ί,���Pe|�-�Zd�_�-�-�GV_� �����d�%$�c�Z����O��?���1��	�x�aI���f(��xEC������I��켳N�U%e�'��s��H��7n\ɪ7p�Iм�0Z�y'��U�	b��LR�<��솬�7��٢=�ؽ%[�e>	�F��EIF�+ɮ�H}���ɂ��)}��J�q�?�f���޵���n}��TsQ�g���]OY�s�[�����;�~�0'Y;�Ǝ�z���F��ޮ^�d�`͑ȟ�ɐ��	��V�߄��m(Qb�G�!�^Nh=�B�HM��mC������ ҥRI�[�1������-�x�AT�)����S�u��Nz����)�%���7!��o�4�te/}v��e�)�$���p��_�������\����"A����o�/�Q!���B> >[	�Aa��jt�vL�"=��$�O��9c�3�؆��<
X�V[[_�J���Q$�B��,�w�@q���G*�E[�\�)?����|��$�~C�% 2�����P�����Tp���%.Ⱦ�}�����=i��;=���g0�HX!/��v%���e� ?���A�"��\�|��G|P༘��Z�c����Lz4d��?2C�%ή��=��8�ܨ�}�ӂN�<�i��tP�nU�=zf��_D�L��Ʃ����F�l�0(fC�j�"���-Ƒ��O�$�F���BLˮ���ͼ��St����P��ya��F�ޥ�P<ƿ襂�ď����I�t�#���ȣ��Q?*⸶O�ȵǴ�� ����G��Z"�ѻڸG3�i��H�A!8T�T���Cv�eTj���I��~�y���AED����)���{��w���,}D��^'�^g,��������u� k�7 z �{^�6^Yk� �Яl��Ђc�����T���y�U(�j.�dB^}s��CR�-_��`A���R,�-S����jк)����P!s��0�✘S�n7��4ڔ'�6f͋�B���$�q��˧_�Ij|_���������uV�yG����èDK�uuSlз�Ţ�)�T1G)�'���"�SZB��O�3�jn�%�(��}�|,�|-�n��q�iB��o޼8�e	MZ���$~�I����,�{�\�t���)f+{�"������e�? �G+�"�{��:�KQ��6�����R��u��ī9=�/���O�(�9��G�N,��d��B���B{�<���9S���)�{W7���]���y&1GQ�Ӥ Vi�3!Ħ��N|��P�x	2͕��#�u��!1f���"w�ݡ:���U�@�/�Oa"�WN3�������˳-g5����G#�m�u@�H:'��l�H��D�BU��c��s��H��_QO�v�.Fp?0&'2^x�3rM �)��z�Wa���v���F��ݻ�¼�TAd�y��0��y��L��͋�D��Ꮏ)+����¢���PS!�5Ϣ�U0|9��a�@�\�ZB}���ح�c:ޔ�zwKsS�~��i0|�_ͱ	�8�z�}GYX��Q��b�mҐ�'����E���`��}��/��H���g����q��E1�tt��tD����RQV s�裂D&���/S��΁�̳%��)�%�#����^���`'1�Z�&�C�y��k|���lِ���~�VVV��bm��tnܼY�����@>��sķwj|�ɤ������a����
Ȩ��� 
���"x�$XW�֖��J�]����HX"�~VH=ca��^u�灑�����q����,.Is�9!�v����)rQ�.��ȸ����>�!ڬ��W\@���Z�:��@*)є����X��-3�ؑJ��C���=W��w�&��dD4��d޵��l����CV���@��!9��&O����ܱ��P�D�����F�p���p$���6ݼy�;�a$�I���(�;+�؁�s�����S/�HII�:ҒyjB"��D����v�ރ�
4c�� ��ȴ�i���`��Db0���ж�X�t�Q	0ӡOyP'(q]&���>=����� u�1<;�Sy��r���K�`F)j�c�lig����A��$E��A�>D�cGM�۷q�1��j��7�`"��G��kE��M#�*x�5����F\�ЫݽGY0睨k���B�Ә��m��|��sI댾uE���Ct����!P\\���<<�:����T�{T���Ⱒ�b�ėtyʷ�v���Ǐ�~8�zo����U$�B.&t.���͌���.P��C���}���|d��7��KUl���\b�[X�m�o��*7�f�wЪ̱����t�cMR|2��>lX;hu�Ru]ר�*ԑ�7|ۀ�i���*�
��?��t�Xe]MϵNSE��=��'9�6���O��%ʼ����G�9��ev��."G�(���~��b�M�=��1�Pp�P��5Th����䝥Rg?F&�q�M�8)�)J�7��7~q��C4]�ܹ��_�$�Բ�k22�D��)��H,y0��
��O����H��/J�*\�R7�5�(�'���[�E�=瘇p��л;�Q_���=܃\#�ۭZwD��x���N�C�ҷ8抱� ����s�{� %C��B�����p��;+\���R��[
�Q/� ϼߖ�)�����^�����.�[|;�iSE7P���`��w}aP��[b0��*#_��+52�YA_y��n!����)�x�'�b�3S�L�E���c(�* J0zw��{:%��t�K��� ��Mx_=�WP�<"�S�m��n��z2�6O�6���P�h�z�K��k�68Xf�3�3w6ũ�
T6��:0���M����C�d�}�7ы��#�ČX`&�b����g�J4����& ��J-ٚ13���*N�FX���+�9��QLsM0 �I����ۛ��w�s�=�DY ���ib�C8�Z��<�.���t�+[b����un����L[��#J\������j�uF�>7ԇ%�_�/����e������Q܆� �_O�wEh����/����y��yE�$@��l TbV��h?����������5����o�O��
�~����G��.D�p4�{�П�9ɼ,I |��@c�&y�uݣc.2�yl��r&�>p/��*..c:zQ ��ẓ�A�+�o��S�x��%$^0�����p�g	 ��\�`�$��1�'<��¸=�{Wl������\��fz*�!�KP�W���~&$�q2$$o�$q! =��P�����O�9���m<ąН?�j���c���4��,��{7��<�_g�֏�F[�YA��g3���p��_��dGGǠ05"�����{����W������rlEE�6�ǌ|�ƫ��?~-C��ٝK��&>*=��������ǭ-�Ԥ���o�r�T�V��!���<��V/���J���S��Nk:���X�OEg���^��n�C�Hv�備|���T����ڪ�Y�A���c���QQ��W9υ����Ӈ1x�0ǘ��._�)ǋR(Dh��L/��� s����j��n������~\�s �<�c}M>Wü3]����T��Svjc}}G�	�Qh�m9{^eV�F$~��I�W�6�v�g�	/�)Fgϛ�������b^����^�����p.,:B�7�b����+�X7{��!h|��
0�P�*8��)����(q�}&�Xl����6�cP���P�?��ZŸ�l�2b�>�r���h�^EYY�aQ�S����w������̬�U�
�&83�:����^b���ݻ�nnn������n�B~����-hk���W��D}�KQY�䭭w'�Ko�|��u/J���Vj��('�^��-̈́��9�n��d;�}lg�w ����$FLKJ-�(�t�ۚ��.��l����̩�Ǝ�%����=aYa�̐�h�l�w�v?z"���ү�#�${Q��D7�3�vh %�����輊�r�jf���1C)��⎿���������c�)�� ���<ُ��)BT+��|��Rת��� �:�C= �ף)'h�5'`�[�[!.�@�aI�J�x�s��U�.��S.��٨;6��K��"����8�}��Q��-Vfƀ���끽!��b�ʱ6~~f��DK�h2J����&Nq������"��<t˱I��LEM�]��(�xnb�H4�c!�i	=��RR�;[���^C��я���4��s��Dw�k�q����ͭ� �_%�p��I$�w�̖ ��bArl���?P�Y�x�yP�?���	ui	�H� ��k3�[o��J��� �.n?;�S�m��[:�Ǻ��y��b|�4xA0���	&�<��:�śWI�U��"
W �$���
\\�[`����GB��]��P �e���g��0C����&�����޴�x\��D�+�kff����-"����P��XM�厹s�Fq�~jI;���9�=�D���d�]�1L+=NRn��#�����K�P�>L@i��I�AN&g�K�hr��"#���E���	�
���L5�C\o(W�V�)id?�VFS�Z�s"�R���"������	CC��30��ւY��!,&h!���F?\�*(]���(�uø���ԕE�l��M�`�[Y�~qJ���3h���<��b�p'�_:h�����\�i�>�����j�������G���٧�����"%| �9��Z�Ԟ��D4W9�À�@��K����%tc��'i����r�GԟV����^?�=uo�fW��|�Gq�b�,�ptu��� G��4�rș�#���j��xC!���J�wd�A��	�Gf��o0������g��ʊ�l����oP�P���PȈᗿέ�
�D�%A-�l�ʚ�T���2��[a�ȠR:N"]ﰯ2��'/��ƛÓn�N�FƗ�HdsKU�CE��������\��ʩF��׵�7�z����<�q(~a��K�
��n�����6L�A.���S�"��a����*�-o�TT�S��ˏY>? �b)�	��\��pQ�<LMOs���9���M��a�~����SÛAfFc}�av������닛#\4̔�F���xw��^.D��X��Ç���1{�;��Qˁ��$|����;	�{锑����>�|.��61���o�����P�GF��M��d�,"O��|�y��w����f���������X:��ߥ�O�;�sz����xU�����=�v�D�u�i/Z<^<Y�ң����|���xjr~�/���ac�����.gl����?3ۛ�Vw�Ly��xvW0��uY�B�3v�K���	�g��h���ĝz�ý����[�r�r.�0ӅgFGG/��Y�8{�}jfV},6J�k3�(�?1c��sza�Z�,}�$C�JG5�Fb ��cT�ԮP!���u-�����P.��œ���E��������]�����m,}W��>N��W��<9A���=̯�g�S��vnw�0���Z�-���@���LML|:��D��;%��ׁ;�( ,Ae�(�p����#YDv����e���1�-��l��N�9���kl���w�z>��6s���|��^�'Q��]�G�k|�nY���>4Lx����[��s�(�r�z�a�e���7��������?����+�YF��A�7U{.~�G��yｼ�(lV3�_�v�t=�o�k�nt���F?�d(?>�-�_k��5�&d������a_��LIN�,1����}0,6��/_��Y��K�n\�Z��}%)3�.���U*6.R��?X��_�<�_jQ�;mS�ّ��_a�B���k����귆i��7nT��h��\{+�_��]*�5;;{�Y)�h�k~Zخ�$���YYO_�Ҡ���;��ϭ2V`g��/}�/rssY����8��ܓj�x��ʣ�`�BAhz����������k��`������r��v�
��w�.^f��n^��?�}_I�䌬,��������(}GY)j�q��?������W�vGq#E瓓�t��F���q��)�>��Y]LL�_%�/ڍ���E�K�e���/�ֺ2}ڴs�ğ={&U}OI��� ��QS���-j�_��j]�6��v`B޸k׮�魁l�u~|z�*+�$�����J��ϻ�m�#����vW�/+�f�4(s����*y�iQNN�����_�� &0/v[\XTW�ov`:#��UW����{�s��;7��{|�w?�7{l�3$U;x���ͮ;܏�� Cp�|��oi1��\hqg�N�q��#=�v�m�Z��j�>c�ϱ;c�n�~�d���V�+Y[+~{��	��ߧm�	,��6A.�j�	㿃��.{����=�{�������j��wr�����~.�� PK   Ci�S�R�η  6     jsons/user_defined.json���n�0�_�j+�`��Jv�H�6ڴWU��ख�Mm�*�x��sP*�d������cs@;�h�ZE�ߒn�%��?*<�s}�Qm��*4y=\��N�&Ίnw�7֌������[��Y~`-W (��n�� ���5;�����9idKm���q��y�qJ������;	)1�c/��5�U�dusJ�ڿd�@�[�-ıB��A5��hr@�ݝ���
C~䒘��]���=�I1>N������6_��F2�BO����f�ġ��cG��I:uuϋ7!!��d��Tϟ-����񁁏���d���<�>=8��� c~��#�jxD�p�5�y��O���~ًOo�,��w��n��P��o�=��ڹ!a���;�|Z�(P�<�"��o�h��[/���/�I��;蒢��a��ݭ�OPK   Ci�St��R$  k            ��    cirkitFile.jsonPK   Ci�S%�$�& �\ /           ��/$  images/66379bcf-d80b-4bdc-b204-78d4e16074e1.pngPK   Ci�S�R�η  6             ��cK jsons/user_defined.jsonPK      �   OM   