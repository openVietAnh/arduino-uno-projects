PK   r��S�QE�  i'    cirkitFile.json��n�V��_��A�Y���'����	07݃�F�
�dIic�F��4�<м�<ӜM:U�h�d��07�Wl�K���6�(�}~�������q�~�;>�fﭸ��c}���>�k��}�{hO������?f����~��7��z�9�}�m�,�m��X��U]l��&�W+[���u��mj����/����tx�=���r�LU��[j��ja���l6�f�-���R���j���?�]<������2@�%DR[��
�-�Q��S�!���:�UHmf�*�vf�*�vf�*�vf�*���E**�),r�(V�#E��m=N�W{z>���O~���2x�O��P���E��=}��ס�o��>��}��CjX"S��a��0L?�Z���H��
�zǏ�E<��%2C�9��i��"E��"F��k�"^;�x�K$?�S�kg��a�Ԗ�������������E�x�,�3,�)�3,�)�3,�)�3,�)�3,�)�3,��*^;��"^;��"^;��"^;�����U�v�%2E�v�%2E�v�%2E�v�%2E�v�%R[�kgX"S�kgX"S�kgX"S�kgX"S�kgX"S _ �kg��a�L��a�L��a�L��a��6����������9��t�aw��w���i?��ǻ�?�Ώ����۠��t�ҥ,�zg�w(��t�-X�
�;��X�Ԗ�w%�Jg,]��w�Jg,]>�`��Y�P:c��ў��a�C錥K��n�z��K��%�ݒ��3�.�+ֻ�Jg,��3
��ɂ�3���v����/�|ap�08a�|����p�`���}a����������i��3���8����g0��+����`>���N,��|~:��>X>����z�3�?X>��|N ��?X>��|6����?
8p�`���$�p�`���/�p�`���Y;�p�`����F�p�`���R�p�`���9^�p�`����i�Mp�`���yu�p�`�����p�`��󹌰�]V�mVp�(��Q����3���������3��g�������3����������3��g������3���I������3��gx��Up�`����p�`���Y��p�`���~ �p�`���N��Lz��?*8Tp�`�����p�`����p�`����p�`���^#�p�`���.)�5�?X>������?X>���3��?X>������?X>�����?X>�����=ۜ�n��5�?X>���w��?X>������?X>���_��?X>�����_���`>�����`>������������e����M�v�l�7q��N��W��,S�.����䗝?'�~ٲs�6'�~�$s���-����Z��kS���];u�����5u����֤���n���ӯ�O_D��/�[��ޢO_��>���5u��go�J����b�������_쓟���'?�`���_?�E�]-V6��̿�?6��?ue�e�Yo^;W�{�ٯ�G�~�s?j���Q�_�ԏ���w��׏��v�~�7j��g{�f[�۪���2ﾪ��zY���M��o��2-���Q�w���n��tho�����O�����K�R���D����딖_G����3Q�_���g� �n�{�J^S"H(y�b� �䕏!���S�J^�"H(y�g� ��]3�J$�ԝ������ S���7�r=����u*�Lϕ��
2a��WB���5���\�:���)��A����ʯ�L��{�?�A&��SJ���V�+�R�p;Ą����R��;�ĝs'��x��qJ�_�b����4�Rꗆ���:^`u�Rꗍ���:^`u�Rꗔ��8V�K��SJ�r�w%��������R�0=Ą����R�h=Ą����R��=Ą��
��R��=Ą��
��R�V����k��Eq��WX��R��=Ą��
�㔒O�Ř�:^au�R�I��W?X��:N)��D�	��5V�)%�D�1q�nr_obu���8���0&���X��|�Ƅ���㔒OH���:�`u����'��p�n��jV����r��
��`5	kj/�5᪠�
V�������
��`5	k�]_/�10(XMσ$�^vi`P���5��H|����8�`5	kj/�9ઠ�
V�������
��`5	kj/�?ઠ�
V���=��`�I\Z�����oE�K�4��4��4�KBkZ��\�&}IhMC���k��$0	�ih�����&�5��a�x�IbZ���\���4&�5��)�x�IdZ�������T&�5����|���eZ���\%���\&�5�Ϲ�x+�FL���&��\Vhr���4�>N�&�IhMC�s�4�jr���4�>'Q�&�IhMC�s+5�jr���4�>GT�&�IhMC�s]5�jr���4�>gWsc�&�IhMC�s�5�jr���4�>�Z�&�IhMC�s�5ފ�Vݮ��e�&���\&�5����x��eZ��z����\&�5��J�x��eZ��z����\&�5����x��eZ��z���&�IhMC�D4�jr���4��E�&�IhMC�]4�jr���4�ޣF�h&�h*�&�U�\Vir���4��3H�&�IhMC뽏4�jr���4���I�&�IhMC뽨4�jr���4��SK�m��eZ��zo0���\&�5��8�x��eZ��z�6���\&�5����x��eZ��z�<���.�6�\VkrY��eZ��z/C���\&�5��d�x��eZ��zoI���\&�5��Ȕx�hr���4���S�&�IhMC�=K5�jr�����N\�J�ۉ*Wz�N]cQ���{�J�y{���D�+��'�\�n=Q�J?�*W:HOT���yꨃ/3z���V|�*s�u�Tf_[�t�3��eB�KO�yŗ��N�z�(.�;U�y_�[;U���V��*Ì�kkAN��F�p��2ϣ�r��2ϣ�r��2�(��=�����k�~�)�f�Z�l�/��\i�lR�,�ʶ�b�ތ8��°�������i�ʛ�Q*o~�F��yH���a�ʛg5�T�<�Y6۲�V�|_�YeU5���X�כf��6�eZ.���T���ϝL{:����i7{�����G8����t\ߟ�M_=J�kE� ��}�"H(u�!��RW�"H(uu!��RW#"H(u�!��RW�"H(u��J}RfJ$W�����m�
7���V�+ޔR�/U0LX�6��SJ����0a5ܰ"N)���Ä����R�/<1L��7w�����R꯯1LX/�:N)���Ä����R�I2LX/�:N)��j)Ǳ:^bu�R�>Cw%�������㔒�����:^bu�R��#V�K��SJ��c��x��qJ��+`LX��:N)�|~���&�]��x��qJ��]cLX��:N)�<_�	��V�)%�W�}�����㔒�cĘ�:^cu�R�ys��&��&V�k��SJ>�	c��x��qJ���`LXo�:N)���	��Vǯ)M��1��C��S& U����5��y>�*諂�$����UA_�&aM���
��`5	k�]_-�&a��A_��&a��(_��&aM���
��`5	kj=hU�W�IXS;�@���*XM���k��&qIhMC��6k��.Q���.�/�$/	�ih�^s����%�5��3��V��$����{�5�jR���4�>�A�&�IhMC�s14�jҘ��4�>�D�&�IhMC�sc4�jR���4�>�G�ł&�IhMC�s�4�jr���4�>�J��1�Wb�\VhrY��eZ���8���\&�5����x��eZ����D���\&�5�ϭ�x��eZ���Q���\&�5��u�x��eZ����]͍I�\&�5��=�x��eZ���j���\&�5���x+�[Qt��&���\Vjr���4�>7_�&�IhMC�=4�jr���4��+A�&�IhMC�=4�jr���4�޻B�&�IhMC�=8$�V�\&�5���x��eZ��zO���\&�5��v�x��eZ��z�����d��d�\VirY��eZ��z� ���\&�5��>�x��eZ��z'���\&�5����x��eZ��zO-���&�IhMC��4�jr���4���L�&�IhMC��4�jr���4��sN�&�IhMC��4ފ�|��|hrY��e�&�IhMC�5�jr���4�ޓQ�&�IhMC�%5�jr���4��#S�m��eZ��z�O���\&�5��,�x��eZG;q��+�n'�\�M;u5zD�J�*W:oOT��+{�ʕ��U�����r���D�+=���:h�2��ڢ�Se��{miթ2�����Tf_[&t�3��-�9U���(��J�Tf_[r�3����8U����5�z�eF���ȔE�]-V6��|���?6��?ue�e�YoF�ՌRaX��@�Ry��4J�͏�(�7?M�T��0�Ry�4J�͏�(�7?I�f[�۪���2���f�^��z����f�L���cw������&���p8�w�g�-��~�;��O���ݶ�{h���8{��×'���D
�s�	<y���Md����J}�"v<�>};*F���ۣ�/��[�|���z|�<��6���zx�}w�>�������!������;����*��W/W�"z�e(�[�"z�e�g���PD��E�@�P���~D�O�t�phO��.�_~?���|{:�Ow����b%��,]�-xE�(�.ϵ1��D�e)����K��ZJ�",��k1A��D��)����K��ZR�",��kQA��D꿡����F��(�E��&HY%�g�/I.��@��4�d5����/H.���P�R� �
R�<����{�@I7���5R��s�(�P�����;�A�����q��F꿶�r '�pv�H��Q��@=�k��օ(PO���5R�D4����i\�ۋą�JPOK���5��#�����qop ���i\�[�@=��z��Vg PO+���5���A\�%�����i\��@=��z���8 PO+���5��
�-POk���5�������qop_�߆���i\ç�@=��z��)� PO���5|j1�����C��Ӂ��9�~�nH�`>��R;�R��!��|�v0m��C�c��K�e�����̗��ߠW���|���ؿAϭ��e�������Z����̗�A-N��3�/��6Y���g0_j��8=�?��`>�]�>��Lh4���I{��<��9�� bt�	�&��di�4M����҉&4���8�=�S	Lh4��M{H'��hB�����N'0�ф~:�!�P`B�	�z�C:���F����j:���F���C:���F���C��+:�tN)�M��]h�M�suh�M��h�M�s�h�M��h�M�s�h�M����B�M�si�M��i�M�s1i��ۻ�R�9��s
Lh4�ρ�=�s
Lh4��ߥ=�s
Lh4��=�=�s
Lh4�ϛ�=�s
Lh4����=�s
Lh4��W�=��M�s�i�M�}h�M�=h�M��h�(�T:�TtN��M�}1h�M�==h�M��Hh�M�Th�M�}``k:���Fz�C:���Fz��C:���Fz� �C:���Fz�#�C:���Fz�&�C|�<>m��)5�Sj:���Fz�,�C:���Fz�/�C:���Fz�2�C:���Fz5�Æ�)0�ф�����)0�ф�׎���)0��E8q%�A�é�j���������|__�r�ܠ����-I'�?h%:q�AЉ�ZwNN������ۦ
��N�����bS��[�뵵��/���*}ӗ�}}�����T��(.R5U :���BM_���� �/������*}1��˯����Ck�*�"P�v�X�|_����6�ؤ:�Xԕm��f�y��d�����C4j�W>C���#4j�W>A���00j�W����ld�����,�mYn�r��˼��j��e���7�~�m˴\�6�F�ߏ��of_������Y�їT�1���0�SR_��?�^"��x)�C�������4��c������n�x���(|����=
ߣ�=
ߣ�=
ߣ�=
ߣ�=�G�c�9�M��Ǹ�E�cv��7�awr?ۼ1�N��.���߲z}$_y,�ӭ�{�?��T=2�T�^ *�D�c_�C�*J:[X�@TG�B�C�DMtlGƑ���-�D�qd/��e�(4�^����D�q��J~��xj�כݽ�N? �yw��W�-��Ɇ���M�pS���n��7U�M��z��y��7-�7-���ϛ��M��M+?�X�߷g��������=����V5e[�;>��?e{�۟|4$?���?�O�,�S���8>펧�]w��ݧ��M~�����÷ف��w��o��}���߾��u[��2�,���??���Yw�~���协�����6���;�������ޟ2f�����~}{z:�?��}�{8 $�����tw�>|��|��o���]�-t���'e�M]�r���4_T�v�N��Xn���E��*����~���ufy3;��{��	fO��n���w-C9��j�>��_���t��Vg[lq��9�R�o)Ϸ��_�g�Z���>�{u�rθ�w��쿛fU�j�lh��Q]�Q}�RZ~�_~���t�Ŗg[lq��>����/�8�%�mY�mX���>�{u��◿�����;���i{w����ؿ��.��\X^�p^�����7o�,{'��M�H�*+�<��?-~5hW;[��n�]]��,�Vٚu1/n++�M��W��A;*O��>��VE����_Fp�j�Y�����q�����W��{����z��,WVcֿ�/[�����W^�ˏ�^D�������Ǖ#��)�����7����g�y{x�R��:�=�sm.R�\���.겗����y�����ۼ��t�����OQ�a��q��L�v��/i2������/��r���������.��+�?��������?�_�����!ep ���w���w������|��=��du��ƨ�(UW�r�xg����GZYV��(n�!�n�����j��������W��vy[�¨��U�;ԅ�.�HϛV�*���1����PK   r��S�QE�  i'            ��    cirkitFile.jsonPK      =   �    