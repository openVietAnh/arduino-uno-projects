PK   "�SKb6��!  �O    cirkitFile.json�ݎ�ȑ�_e��US����n,� �5l�c�F��"i7��K[�������3m�%U�T����.$u���`2��dF�x�[��h7�]����=�mn^�����j���:����y��>mۿ�V��z��G��x����X��U���6mW���uW��鋘��hVkW4�TM�^�u�Z׺��o��~���\+fU0�7����_����`f�*�6��
�Mf��kK3�U����������`Upmcf�*�gϳf�L�2On�߿�>�O��k�P�+�"VRM(�EYu���wq��oLIR���ژ�ś��m�bܽ؂��g��z��~�h:����v��>�v_Z��m��co���%2���j�p�
����/�f	���y�m��z��1Kd
���o�Ҙ%2�݊�%2�݌�%��~3�=w��4|��v�=��K�S�Y��P�Lј.��x9����o�w�nuw?_�}��_���Q<���vM��%$�/!f�La����J֞�f�����,�)��D��_~���>t7Kd
���,�)����k�}�n����k����k����i��������,�)��,�)��,�)��,�)��,��dϝf�Laϝf�Laϝf�Laϝf�Laϝf�Lxkϝɞ;��;��;��;��-��,�)��,�)�s"��f������G�탗wL$zW�@M$2�	Ln��lq$�9;�`�K�Z�����J'X:�l�6vP:��e炍]��J'X�<r��.ac�,]c`cWbc�,�k+l�*l�t��sm��]���N�t�m��k����	�N_���cw�	�O_S��.���/l0�0�|��W����,����5mp��N�'`>}�?����	�O_��8�|�ӗ����,�����|p����'`>�X ��}`�̧S"�7����'`>����`�̧�P��C?�@?� ���?�|�ө?�����O�|:i	?����	�O�[���X>��lp����'`>����`�̧�����,���^N̓��q�,�,�/x+l_�_�.�}	`���0�N��l_�|��	����_�B���/l_ؾ`�̧�^���,���t�.8~`���0�N4�l_�|��)������O�|:�?�}��	�O��c���O�|��	������O�|Z
 ?����	�O����X>�i�p��E�3E��#��G�,�����8~`���0�� ��?�|��2#�����O�|Z ?����	�OK�`����'`>-J��`�̧�t���,����8~`���0��0��?�|���K���'��g���G���X>�i�+p����'`>-���`�̧E����,����<6~%�`�̧�����,����$8~`���+|���%\�̘��q%��͏˟.��g[R�(H�D{���~���ǅG6?����q�ϥ��z2�1��%���?.仴�q	ޥ퍝o�R��#����ԓƺ{oٽw��G���k2'����d��$پ��j��Wѱ�>��^iڽ�|�JcƮo�;�z���3���RXK۟��_vM�H1�!�w���K��*E�j�^�/��g57��|ڙ��|֙���V����Y��_�g5?�����XsV��c���^�/�����k/UQ%�m\�>ȅ^7���^7���^7���^��Z�2�b�
�"�n(겔bӔ}�R�1��}V���}V���}V���}�tCS�1E����d��}L��w����q���K}ʍ)b7źYu��J6Ð�ns���i~~�]U�1�$��R�W��up�!U������g5���ؾ}ڶ���vw��G˕+����X����/�!�ʯk_�1�u�"	9=1D !��QH��Crz����� 0D !�cH��0Cr�]:P��e�}��&��Z�L�ҷ�6������J�$�Lϙ[���K�{%��M�sn�64F�Q��߸7�62�Y�I΅��L����ͯ��	��QJn��b��p�%q��o-��`y���8Jɍ7�AL %7ޙ1�F���QJn��b���=l�Rr�v,����[%3,�{XG)��V=��Y��o����P�.��x��q���u�1�Jo|����Ȅ������QJZ������QJZz�����QJZ"��G�x���<`L�<ay��%'`L�{⸛�<ay���`L�<ay����aL�<ay��ӷa�~`y<��8JI�Ø`y<��8JI��pO7q�7ay<��8JI�B`y<��8JI����`y���q��N-�1��x	�����q��P�q�ש�n˧�MY������D���X��*V��P����`
�k�+��U�qe�
�5�.J\��`"�`
kQ�z\o�PX����:,�0X������,pU`\�Bau�q��*0�V������\W�PX��`�1`���
�V�m�Ė�H��㻄c���(�¡�w�9��/
�ph��yNl9�B+Z}��[���
�V�0pb�qbZ���\Nl9n�B+Z�S-ǑQh�C�sc8��2
�phu���ǗQh�C�s�8���2
�phu�'��'b�Gb_�9��s|�V8�:�[�/��
�V��qb��eZ���DNl9��B+Z�[ɉ-ǗQh�C�sD9���2
�phu�+'�_F����弘�yC�B+�iA�����eZ���jNl9��B+Z�Ή-�mE��_8�,p|�V8�:7�[�/��
�Vkpb��eZ��j�Nl9��B+Z����-ǗQh�C��+8���2
�ph�%���B+Z�%-ǗQh�C�5Q8���2
�ph��'�_F��֨�Ė4��4����"ǗE�/��
�Vkqb��eZ��j�#Nl9��B+Z��ĉ-ǗQh�C���8���2
�ph��%����(�¡��`��r|�V8�Z�[�/��
�Vk�qb��eZ��j�9Nl9��B+Z��ǉ-����Ǘ%�/K_F���2�Ė��(�¡՚���r|�V8�Z[�[�/��
�VkdRb[r|�V8�Z�[�/��
�Vk�rb��eZ�G�y��U��.ơWvE��.�P����BYI��ϭüP�Lmڅ*g��.T9S�{��s���w�������l���n�P�L=�*g*H/T9S�yi�u^L�L�=���R�3��ʜ���TӅϭ9�T�ޟ��K/�y��ǫ�.�zc/�.��T��[�TӋϭR�T�/��Tf����ߖʌ�x���R��^|�~�R��^|�\�R�}/��Ľ������V�,|�5U#���<V��_k��_U���~�Z���R��\=�f�\=�f�\�(�R�zM��r��0K��a���Q�,������S $_4}_1�+�^��J�۸�W}��}w��վ;K�jߝ�r��6����جª����,��4e����!]��,��q��r5.�T��e�tCS�1E��-�e��}L�z\f�\�/U?t�O�� E��X7����\�fR�mf��9*WY���c�W�M�B�˥+����B�&J���u�Y*�,?�2�Ӷ}|Z=�7��,�|�{�?<�V��|�Wa	��B�@Bn<� D !7��"����"���"���"���-"���@"���S"����q¤H\�ƥmX�X�F)���5,w,y������	����QJn3���K�(%��M�a��q��(%����a�qpX��<�Rr���&X��<�Rr�;�&X��<�Rr�{�&X��<�Rr��;����QJZ�Ƅ���������QJZW	�����QJZ������QJZ7�����QJZ������QJZƄ�'��)����QJZ� �����QJ:_�����QJ:?����,���t>0�	��,���t�)�	�t�x��,���t� �	��,���t^�	��KXG)�<(,���<~Ni���ɜ9��~�@U(�Bau�d�ZW�PX];�+�Vƕ�*V�NꗠU�qe�
�5�.J\'�K `�
�5��(q��-�D��*�<F��uR��PX];�W�Vƕ�*V�Nj��U�qe�
�յ�:%hU`\�Ba�w�9ƀ�(�¡�w�9�%�.����.�/�8/
�ph�]sNl9�B+Z}g�[���
�V���Ė��(�¡�9��r��V8�:�[���
�V�pb�qdZ����Nl9��B+Z���y���eZ���\%Nl9��B+Z�sŉ-��Ǘy�/�_F��΁�Ė��(�¡չ|��r|�V8�:'�[�/��
�V�Vrb��eZ���QNl9��B+Z��ʉ-ǗQh�C�sv9/&q|�V8�:��[�/��
�V�Psb��eZ���\pNlIo+�^W�����e���(�¡չ���r|�V8�Zc�[�/��
�Vk%pb��eZ��j�Nl9��B+Z�]��-ǗQh�C�58(��_F����Ė��(�¡՚(��r|�V8�Zۅ[�/��
�Vk�pbK�IF�J��e���"ǗQh�C�5�8���2
�ph��'�_F���p�Ė��(�¡�ZT��r|�V8�ZS����eZ��jm0Nl9��B+Z�qƉ-ǗQh�C���8���2
�ph��'�_F�����ĖT�T���Ǘ%�/��
�Vkrb��eZ��jMFNl9��B+Z�-ɉ-ǗQh�C�52)�-9��B+Z��ɉ-ǗQh�C�5K9���2
�̣��T���k�P�+�"VRM(�EYu���wq���a^�r�6�B�3�d����P�L��*gje/T9S�z�ʙz�U�T�^�r����^꼘�{n�ץ2��{niե2�|nӥ2�>|n�Х2�^|n1Υ2�����V�\*����ւ\*����V\\*�����5\z����s�~�	�욪�b�C+u���K��*E�j�^�g�jf�`X��P�T��O�T��N�T��M�T��L�T��K�T��J�T��I�˧@H�h��.bW��TE�|�q��� ���,��}w��վ;K�j�mb-U|�Y�UC7uYJ�i�>V)�����R��Y*W�2K�j\־�H74E�PD����YPVM����e����R�C����R�:n�u��
ʕl�!��fFߝ�r����>�|�t)d�\��.�/��j�4~]^g��r���m��ߟ���~�kﺿ߼�p{��ݮl�߯6}��=��]��n^�}�y��iq&���ְs-�y����@k��F4��{۸̺�h]Zw�lcdk�{1_l�^�]O���x������/N[�{�G7��hE��Bo?� ���fG�5�EŬ�)8�5Aj��-����n޽�8f���o��-������m����_�����9�0@ƾ�X���
�HCac(��bL���1�Q2��:X�PX��?w��?���z�9y��y�5(Қ����݂��s�5��6���A���wf'��q�w���a�>>����ן~��^�}ڶ�?�R���:�6J�񶾑B%��?b�v(���J)�n|Rm�0K��I���,��'�F
����)�n|Ro�0K��I���,���?Z�"��H�ވuB�4R���u�xB�2R�度�4���IF#�	��H����HyB�1R�]��ߦ�r R� r�]����r Һ�u��ۿQl�0k��+�V���R�]��_��r �0:�k��k�V@>��>��.����bҫ]��_4�r4��F�n��:��@���k�Е �a�톭.� ��� ��v-�� �� ��v-�� $� H�v-� �m#`lk��"� @z���j���� �m_�}_@>��|j��� @>��|j��¥ @>��|j�Ђ��'�|� �Ԯ���|� �Ԯ�� �i�'i�|� �Ԯ�E� �|� �Ԯ�Ź �|Z�]C�>8 ���ө�������V:z�c��)�)2�5FwR
��0���\;)��Ӄ��'`>�NJ-�� ���	�/�p�&u����'`�<� �oR+��}�|�ˣp�&�����'`>�NJ�� ���	�ϵ���8=H��|�s�1N?,����EL� ;�4��	�%Rt�.nC�>D�FD�NL(hB}C�
�P�F��H���&�w��1D�0��	�Mkt��L(hB}KC�;
�P�pG��P���&Է��1D�0��	uf�F5ڧ�	M��"�1D�0��	uF:��'&�G&h���>ţ}
�PЄ:�C�O
�Pg�c��)`BA�&t�>L(hB�}��!ڧ�	M�S��1D�0��	u�:�h�&4�˪S�B����r���Ё�-S`kж%�m�PЄ:C�m
�P'n�c���ڶ�m	h�&4�N�E�m[���&�ɾ��m�PЄ:QC�m
�P'Y�c��-`BA�qtѶL(hB���aD?^
�P'�c��)`BAjQt�>L(hB-���!ڧ�	M���1�OL��LA����)�S���&�"��}
�PЄZ C�O
�P���c��)`BAj�t�>L(hB-�aB�0��	��:�h�&4��A��S���&�BC��}
�PЄZ$	C�O
�P<�c�D�E��)	�Sڧ�	M����1D�0��	�(:�h�&4�4C��S���&�bl��h�&4��C��S���&�"x��}
�P�.\crRq�������O
�.^��rE���^��PnR�ta�I҅�'�C����\ڻ����?��A���-���]*0)λT���K�-���iiћ.V�ru���_^0o��󗗶[�g���ű���|yy��k#_^�f�^9�x��MW�z�*�R�g����8,�c���R��:��k�F��yd���.忪���z��8���޺��ج�ΰY�/\&f��p�����EbV�׈Y�/�Uf��0V\��!������Q\��RU��ƕ��É������f����f�����XKU_lVaU��E]�Rl���UJ1�t���j���j���j���}��nh�:���~�)�}������)\����_:�U?t�O�� E��X7����\�fR�m.��9�/쿫�>Ɯ�7]
ٙ������i��(�_���?��~�?��|nw׵O�6f���͜����7j�tҠ^����]���Qy:0��������Hd>�~X�Ӣ��h�^[�Q[[xmᵅ�^[xmᵅ�A[�Kۻ���$4?�9�������d�9��sCE���^4��S���a�I�'�#mޘe&���S���U�M#�)Q�����	�h%2�n�D�Jd��'�J�����:j���ҏ�TϮ�D�~�N5V"S?�D���;���GO1�pb�i�XO����޿���6.sl<.H`��;���v�׆6�9�ٮ��Ǧ{O#����O��j��� ��dRS���+��Ѧ�)L7��Mq�)=oJ�M��r��z�TM7�ϛ���yS3��7��&y�$�M�L�ɧf'�}��L�(Ø�������=�wö��{|��2�k����v��Oh���i��%?���߬�VY���W�m�����~�<߿��������{���a����[oo�����?}=�=��2�M���_�?���Mֽy=����������n}��ݮ��w���y��1s�_=|V���~w	��c$�����@�Qrν{���8�-�ԯ�t[��U�!T���F�[��mB6/����+��E��7U�bԞ�}���a�o3�M��lww���7��_m�v�����e(��mj��6�����`K�.?T�[��-�pK8��~�>U�>�>�26�*6n�&�?T��P�k�Z�O[��=~�Aʃ����Hu�%n���~p[������������߿���=}��������=���r�$'�'�q��G>��ϡ�oc�^E�1w��o�l�K�٬��O��jirdV��(aU�!5��>;�>����W͋����Ʀ���������(���<um[7���Q�?���(����6�˝��t�?0�����=�g>�	%�_�c��?��2��~�����~�O��������e�����7�ӕ=�2�Ac��b������K�|��]>��Q��n������B�n��8����	���nx1B���B���ل�r'?7���7�{c���2퍍�3κ;�3� �Š�dW��}'_�ކ�.V�l~�S�/����A9�����O���C���w��Q���::�zH��������/��[w�dk��>�k�˃v�u����c��mx����S�{d����z�Ǜԯ��������?������G�+�'���|�݇�����_�z��=^�;����x�G@��4މ��+x^�^�}G�h:� ��D�7���X�V�p1�)�R�Kb�6�&M�8��1�����r���ۏ����.����Jut%���𕋢C��j�˱v�Yϻfu��aD����`��+ɗ��_����.]_���ɶ%Y��ǰ����Ф<ُO}���O�PK   "�SKb6��!  �O            ��    cirkitFile.jsonPK      =   �!    