PK   ���S��U��  �[     cirkitFile.json�\ێ�6��B}�rH�Ҿ�� ��@ۼ,A��D�W��r�"迗��]�m����!Yk8�����/IW}4m��v��h�]�m�;N��Cխ>U�O�,ylڲߖ���Cr��}O�?M��><n[���b�~8K!���X��km�5�2/�&W�)Yrw?�l�\Y�k]�T:�:�x�Y�e]/�Z���d1�۪9��!�	Q] ��9�h^I]���N�JՖY-ӂ	�Jc�`+��f`�;a�c��2�
�<C,׈�3<���(�A�s�<� ?[��� �8?�@��nA��?�G �����Ρ}R] �}�\Xl �5�_k��O�<t� վ:-�j_�F վ:�3 ��n-���Ղ���j`8�4l>��2�}n)0MD֦�/&ǈj�_<@T��0~����!���şOg3��fہg3ɷ��Wߩ:fI�-�+��;@
l�JJ@�pR޼)�~=-%�$���>�E
E�"�H��L+��@��bKv��ވ���ؒG�R�A]$��A/�_�\��<�#&�y�8(�8(�H>8�)�)�)�);l��#D�ů��3��x�X� t@1g,�Ȯ��&�C���)�D�� �&��g;4O��Д;���\M�	x)�Vl�S_��C���q}p�{=��[�g<�9h�i��g�1Ĩ���9���Uo�$�5���6`��K�(R�-)�I&.��'���8�"�HQQ�dQ��(R�(R�8���8��q������0��`�<�y�8(�8(�H>8�)�)�)�)�)�)�)�E��(N2q)ql�����L\����d�Rn.��$�rs)'�P	�q�{;�	O2#��೨�&�����e����q6K>5�ٕ��jiV�MB���t��=���3��B��c>�Tg��ET#�5�:�R>Ձ^9�@4{VV��/��8	R�9�}�e���u�a��z��]M9�{k���N;f��"X ����� ��c�j���q@7��z��Nӹͪ[���*��}�^'O%�}�B���L�C�Hcq\˸���E�,g ���_���Sh�b �dcs<�8��������.�(>9
P�"tH�!((��$ �!G��Q$�D�=%�DB�H(	E"M�G��.�A/��cy��q�X�b�bq��冰���;� ��JDZ�K��_Y}�e�b�!���ZC2牥�v9�t�te��yѵ�&�N	@�<6C�\��YN�r��U�s	fH��.{9��܈[��]��8f�%�.�p�t`r p�6$�C~�]S��rט���5�=w�q��A�� �A���pf5�'x�A�pb�52���w����aoM�F�<ܿ��(�4Voصi�d4�s���Xi�ea�����xǀ�,c�������������V���jaE��Ƌ��V�o��/�A����w��MU����6����q}���#��It$ј$�$1&�#I�I�HRcRv$ec�>����I��TI�!�ͦ�;S��mչ"�z[n�]�NT����vv
�JQTi���6ʖ�d�X��L�T�����2�yq���Ƭ{���I�{U��}�ex�S�}4]ߘ!�yxl���]�5�{۳�zp�u�|�6{�M�¾m���������c���L���fg,qg�wͮ�7��Yg~�7�Y%w�����ݯ�e��LwM�i�g+^��u�o�o�oW{�c;�[�?lwM?�⽔r.X�u~Dl6+��+*D���v����[		;����ZEʖZ�b��4�Yn�L�j��"��]x�b�Y��l��`X����M�ܘ���L�Ռs��{�h�+�2zz"�91͉v�'���X��#�b��[����W���ן�L��͹�4��ê��:���&%���NfVd|N�y��g��ZI&R�K�d˴bT[��D+-%]'(��N׼�Џ��
��SH��S�b����=�?!i:#�R�}$n���Ư��s>:�I��+��/�2�it�O\�S|ngy���`�ع�Ɂ����(B�(�˓yyt��f�����s���DI�o즧�H���ir�����=����H��?�R��-��{o�N����]�6�?��#�{�y���W�zWar&�*R����,g�r-��d"�MUU�p�p�]��:�e��䥭�Y�L����#�p�uw�����f�y��0i�|�ӶYv�����"��"hG����T���O5���T�Q�o-�şPK   ���S��U��  �[             ��    cirkitFile.jsonPK      =   �    