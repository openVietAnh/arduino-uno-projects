PK   �S����*  ��    cirkitFile.json��n�8��o����K�V��O��3����)(Q�66ˮu:�{P����k��qV�}��U|�w�ˍBg:e��
���!�y�;,������������d���)?��������|w{wx�?��!����߷������a�e��6[���l�b�S�.|t�fe��4M��z�}���o��|4lA�-��~���������6Y/E��r9e�J4*��ͺ���|�t3�O��fX�Q�`�4�5���nX�Q��G44zPC?��5��qHC�0�aG-��4���p���ʰ	��V��V���X�M0�P�bܨ��}�w.�&�b�{�:��/4���`��.&��8���x'3lB�A߈�qT��~ƌ�3�&t���8��@�H`��3�ό�0f��1��̰	�z�a����&t�R���ތ��a�=!��1ێ��aL14i�S���aL1�h�S���aL1;�M0�x�6��s�S���aL1;�M����&�b<v�`���9l�)�c�	� �<��n<v�`���9l�)�c�	����&�b<v��?;�M0�x�6��s�S���aL1;�M0�x�6��s�S���aL1;�M0�x�6�a<v�`���9l�)�c癉����>��|��{��������߹�G�������KGX:�O�~�;gz�d��ٕ��!t7X�5X�t������b�������v����t<��j��A�K�#�v����t���E�vP:���C�j���A�K�V�	����tm�'V<g%X>���`���:� �N0�a`�������gX>�Y�`������|m~4X?p���#0_����q`���敃�gX>�Y�`������|m>>X?p���#0_[ ~��?�|�k�����,���*
�~�/�O��À��?�|�k�O����,��ں�~���G`����8������U��?�|�k������,����0�~���G`���<I�`�������X>�Մ`������|m$X?�,+�4+p�a����X>󵵧`������|m�,X?p���#0_[���`���V*���X>�5�`������|mu8V?�?�|�k������,��ڊ|�~���G`�VK �8�����UA �^�^��?8�p���G`�Vy�8������� ��?�|�k�>����,��Z��~���G`�Va���X>��0`������|��X?p���#0_����`���*	���X>�H`�Ы���������`����N���X>�Y`������|��X?p���#0_�R��/��,��Z}5�~���G`�V�8��������N���6��� ���UHw6?-���i�ϝ�Ov�l~Zisg���;��ֶ��6�n7�wg���m?�yg���m?�{g���/���|��{ҥ���(?gܑ�O�g�#g?n�5rv?tv<{:�<�4tv;�uCnwܭj��c~�GO?�xa��c�GO?�z�ό��h�3C�w����#�%����Ӌr�8��b��ݚ�jηm���������MA�V��zy1*�Z�U���l����峓[��ìg��2�<�Q9���뢳/g�j~���d�N^+
�w�q�Ln]h�u	�o�����{��u�ZbdO��7j���u�j"�q����]�S��J�ssW�mL��%7�v���ٻ�_>���֧E��9���Jk��;gm����>k�:ϊ�,�M�j
qR��u�m�Ѧ-��i�q�z����'���8^��q�*���P]��k�i������������Ԥ�Q+߽�P�!,[O\O����Z�e�ıZs��W��>�s�qb��-��i�qߋM5�ּ2<U�..YU�ͯvn�z޻�_>{	����Ņ��Q2��]��
wb�B�8{W��gO���8R��L|�8X�`�*�3Em\�|����[���I��r�v�(��d�B�e���z'�����M��YJVQ��E&~n檝ZW!x*�n�|W�k�e�nm=D��wo���M�m�����w5߸�����0��rA�����RkZ��Λ�����ג��o�2��%��W:��Z����j��ǭK�:��L�'乛XV��[c������q���d�����u���&b�Y��v[=lW��g�JLquLۢ�ӵ�Ĳ�Hd(R�S�8{W�8�VcL�������w��_G�R���[g�j���բ��I�u&�ģ���=�K\�Z]�[}\O�Q%��PbP�x(��)�I��xPT۸ekl���x��������������G�#&��/����w?���6DZ�8FD("��d���cC��N�#�("��d��ml�~�~�k#�(���d��eC���6cDE�P��7�GC�v#�`�Q��o�[H�Z�_2��6�7���U��l����(K�w�GK�d��o�p���ǅ�����o3����(Kǯ GK�w��L�8n`qe����-�_'~;Ȅ��8n>G�_�~4�X7�8����oAL�8n`qeI?�`q���8ʒ>~1�⸅�q�%}��b��q��(K�|�	�-,��,�2s0&X��8���ʡ��`q���8�R+�c��q��(K���	�,��,�2H0&�;q�KqXw�8���J���`q���8�R+�c��q��(K���	e���1�⸇�q��VN����Q�Z�,�{XGYj��aL�8�aqe�-#�1��x��q��������/Yڿ��t<��q-2�*�����R��d�U���`�@]OW�íu�`%V}8���
�U��DX9�����F	Va�q����5�0
H��+�QDt=��Q@��DX��Z�*PW	VaՇ�*bp�@]%XI�UN����u�`%�6'XDX�ɸDhI���m��V(�J�d�.�I�H&��%�6�\F[��K��dhۜyme20Z��ms�e����DhI���a��V&�%ڶCF[�lL��dhۚme22Z��mkcd����DhI������ ���Вm[�$��L^&BK2�m͕��B_Ą>���eF&/32y�-�ж5p2���e"�$C����h+���Вm[�(��L^&BK2�mm���2y�-�ж5�2���e"�$C�ֺ�h+���Вm[�+31I&/�%ڶ�XF[��L��dh�jme�2Z��mk�e���(4]Q&/�2y����DhI���͗�V&/�%�Vc@F[��L��dh[�me�2Z��m5d����DhI��ծ��V&/�%�V�CD['���Вm�%"��L^&BK2��&���2y�-�ж�.2���e"�$C�j��h+��Lh)�L^�d�2'���Вm�$��L^&BK2������2y�-�жN2���e"�$C�jQ�h+���Вm��%�����DhI�����V&/�%�V�LF[��L��dh[�6me�2Z��m5�d����DhI���Γ�V�ʇP������e^&/�%�V�PF[��L��dh[MFme�2Z��m�%e����DhI�����6��e"�$C�j}�h+���Вm�Y*��L^&BK}�?���6Y/E��r9e�J4*��ͺ���|i�V.Ԧ�i�B5ٝV.���i�B��V.���i�Bu�V.ԣ�i�B�V.�|��u ��x�M_����省U���x�L�������''>�3~����o��7�=y����{�Г6��s�5�ًO���k�����;�5�.�t��f.����ы���s����O���k����[��5�9��L������K�>3����UuzQ.��T��Ú�[�^����X�ʲ�~�n
*���-/F�P�j3��,]V���[��ìg��2�<�Q9���뢳/�Y��\eY&K�~E��V�5��ɭM�.���,]V��x��\砪%�O�o�7j���u�j"{����U�蒟T2����^gbV.�i�s�X:X��\e����O��ձb��%x���-�I��_��\�bMQ�Y�e��^M!N*ټ.��9����X���^��4�ټ�E�0�gǹXY]L��2u��c��3={WL�vE1:5�d�ʷ�.TjK�3�c��sd}��-��sT��{^u�?��ǉ��:��+����T�j�+_UV7.YUV֯vn�/]V����KY��\����S�SJ�S�ľR�Y��\eI���8@��L|�9b�`�*�3Em\:��.+WY�v���d�'q�(��,v�B�e���x��e�*�)v6K�*�{�ď�\�S뺦���uY���.Kuk��r�+��=GO�&�6[Z��/]V��K���*L|]Фr>��ԚV���r���<M|��Ѷp�.Qe���/�В��q���\��%V��&�#2�ܫ-�Vƭ1�Ɇ�t�n����Qe��.+o_��Lm:���h�1f�r�e*1���%���t-*��*�Tx�X��tY����xDfb�a�½=D�I)�Z���.+���Z�XLj�3q�&F��i^���j��{�\{s\%5�(���|1)�I��x\X�`�c\�e�9�G3��������޼��'���(k|w�Ǉ��9���@��rAȐ>�-����wȐ>�Ň���Ȑ>~]����
Ȑ>~�����Ȑ~��	����۰�M������>:a�`��`�eI?}�0��7�8ʒ~�P�a��p�q�%��	����Q����Mn����⸁�q�%������Q����e,�XGY�O߽1L�8n`qeI?}�Ǥ�8naqe�ղ�1�ޤ�^��⸅�q��Vs����Q�Z�;,�[XGYj5�`L�8�`qe����1�⸃�q��V3
Ƅ{'�{)���Q�Zm,�;XGYj�d`L�8�`qe��.�}���q��(K�V�	�=,��,��0&��M��MX��8�����Ø`q���8�R[�c��� ��(Km�0�	�,�_�����zr�էe� �$�J"��p��m��+�����:r�U���$ªg���V��J��+�]"�����( �J"�<����D	Va�1���g� 
H���>���B[�*�J"��pV�m��+����Y/�U���$����$2�-�ж��2�
e]Bi�L�E2��d^"�$C���h+�}�Вm�3/��L&BK2�m�2Y�-�ж52��db"�$C��b�h+���Вm[S"��LF&BK2�mm���2Y�-�ж5>2d�2Z��mk�d����DhI������V苘�'1�����eF&/�%ڶNF[��L��dh�Z>me�2Z��mke����DhI������V&/�%ڶFTF[��L��dh�ZWme�2Z��mkve&&��e"�$C���h+���Вm[C-��L^&BK2�m-���B���+��eV&/�2y�-�ж��2���e"�$C�j�h+���Вm�� ��L^&BK2��惌�2y�-�ж�2���e"�$C�jp�h�d�2Z��m�Dd����DhI���D��V&/�%�V�EF[��L��dh[�m�V�	-%��˜L^�d�2Z��m5�d����DhI���>��V&/�%�V�IF[��L��dh[-*me�2Z��m5�D��2y�-�ж�`2���e"�$C�j��h+���Вm��&��L^&BK2��朌�2y�-�ж�y2�
U�*�!��y�����e"�$C�j�h+���Вm��(��L^&BK2������2y�-�ж�"���L��dh[�Ome�2Z��m5Ke����Dh��������&륨�W.��R�F��Y����/�ü�ʅڴ;�\�&��ʅ:�;�\����ʅZ�;�\�n��ʅz�;�\� ��ʅ��{��ｴ��^3�����^3����^3��M�^3/���^3����K�T�5���K{A�5���K;.�5���K���u1^|i��gf���R��N/���T��QsXStkҫ���+WY����MA�6���Ũj]W�c&s����Ur�Z}����\Yf��9*gt�z]t��:K���,�d�N^+
ķ�����Ln]h�u	�_g�r����:U-�ux
|��Q�}��T��,]V��D������l�U�:�r�M��#����e�*��Wd}Z�����_.���o�s&P��tY��Ś�γ""�^���B�T�y]fs���9�r]���iv�y�+��a*ώs�����e�Х���gz����-�btj�ɨ�ow]����g�������j�[��稚�����7~���{u<G=V��K��fԚW�"��n\����_���_��\e)!�����0�3h9p�֧�j�}���tY�ʒb5�q���Ns���:U�g�.ڸt<G]V��X��1R��rO�|Q�Y�2���49������US�l��U�3���ɹj��uM�S	��9�r]]���֡��Wķ{���M�m���_��\���s��U�����I�|�q�5�<*�=��c�*K-y��^+�m��]��.z��_J�%���uY��O�K�:��M�Gd�W[V��[c������.+����.�]V��"�92��t.<X-uѮc��e�*�Tb���Kh���ZTbeU$2��ر^g�r�?Z�1&������ƅ{{�D�R���,]V��ӵh�cRk���7��0��LO���VWcG?�c��؛�b(1��G�<n�I9L������k�.+�Y~x��+7��p�p�-�yO���_n֏��>���������7��z���+���߼{��/5{5xv;��j��~�������i����+�Q�q;c�O?�w��~�����</�~�����͐�G<3�z���OzX���3wJ����?}͠��o�����۟�?��Z_!�ۏ]!�CX��H1:��@��k1�9:��P��r1��]��C1:�P��1�aƸ�~���?||̏���/?���d��x�t[n�?�^7����j~����|��4E�Pf\�a�8g�D3eǡܸ4�&�q
�4vʏC�qi�M���i�T�J�����	�'��1�	 qx܆~�p{�N��b��q�i��<q�	��m�)�'�A,@H&@L����H��3b�2���4i�d�� �� B��4��D��A�A���d@h6硙�� 4���O��G9 �� b��4��| ����OkF9 �������a�^- ���h[_ 8 ���鸍���O- ���h���xj�t�F+� �S���6Ziq  �:@<��JV8or�r���鸍V6���O�m�r� @<u�x:n��9���J�8 ���鸍Vj���O�m�� @<��x:n���p ���q���O ���h�� �x �����i�g��p���c�#0��Φ��}��0�9�pq� r�Um�ك��#0�>�U��ك��#0�`���a^/���|<� �wV�z�z�|��aX���փ׋�#0�>�U��ك��#0�>�U��ك��#0�>�U��ك��#0_�	��		��Єmn'ZCxOC�y�Bg"`BB�I�h����Єm�/ZCtF&$4a�������		MئV�5Dg&`BB�i�h��	��Єm;ZCt�&$4a������		M��_T��0!�	�B���<LHh¶*�!��	��	:O1�<Š�0!�	�����<LHh¶t�!:O��-;Bk��S���&lK����0!�	�r/���<LHh¶T�!:O��-�COA�)`BB�%�h�y
��Єmy#ZCt�&$4a[���>�>���Xt�b�y
��ЄmI,ZCt�&$4a[΋����		Mؖ"�5D�)`BB�e�h�y
��Єm	8ZCt�&$4a[��С�0!�	��{���<LHh�V6 �!:O���<@k��S���&l���W��������S:O����@k��S���&l%>���0!�	[y���<LHh�VZ�!:O����k��y
��Є��ZCt�&$4a+ǃ����		M�J	�5D�)`BB�2Hh�y
��Є��ZC��y��yt���y�G�)`BB��Yh�y
��Є��ZCt�&$4a+Y�����		M�ʭ�5�<LHh�V*�!:O����Ck��S��t�p�>�g%�n�;�������g�Vw�?+����Yiӝ��J��lVJtg���;۟����?�8�����50��[��50�绒���|�4���Ƿwrݿ���������3t����m�ߨ{{w��[no������o���c������ۿ5���t�7����m�v�ۻ���G����G�,!ťxU�^��ũ4�氦�֤W�ʆ�;�o���l�T�+�Z�Z^�ʡ�u�>f2[��j�q~r�Z}����\Yf��9*gt�z]t�e��]�7οL��䵢@|������օ�Z�P�����o��3�sP�S{
|�Q�}��T٭�w��8t�OaJ*��]e�11+��4�9R,���j�q����O���q{bO�%x���w�ڼ�]��?�u�Y����⤒��2ۘ�M����~���j��a��#q ɳ�D��.&Cu�6������7{WL���S�NF�|�B���l>=����j�[��'����̷s����m�O���_l�Y�����~qɪ�v~�sp�����~��%�R�f~j,���"y�v*�EW
a��]�7Οb5�q����q���:U�g�.ڸl�W���[��K��r�v�(��,g�B�e���L��o��;��d���g�h�کu]S�T������[ׯ�R�ں�\��o�=)�H�li5n���j�u��ϭ�Ta��&���ǥִrߞ��O���ג���2���%��W:��Z�7��j����K�:��L��/��XV��[c��������[��d�����u���Ԧd�!\��v��oW���O%��:n���ZTb�T$2���n����V�_�1&�����Ņ�O�ΣI)�Z����w����ji�ZRk���'��)�HFO���VW�f���~k��Q*���c7�2z�aR%%9�6���t�:��n~jw[��6�����7=i����oZ��R��N�W-�o�xK�[���ԖZ��cw̼��.�_����~���Sk@��i-��vkaZ�Z��´��0��i-lk���7�nz����AO��AO��AO^�A�@�E�����=C�*u�m_��c0�R֎��K�:�{/��c|��Aπ�E��Ћ=C�z�/��1(xy���=��Ko��'_�RG���AOO�җ:������_������OOq�n}la����ɻ�c(x�=�M��+�9��ۿ��Л��
�y�]�9�z��_r�@C/�� ?4�vۼF�z�}�}�(�}�q��Q�!���M�DC�ΉH�~�9'�fȳ_��4�͐gOϻ������y^?���ĻZR����Z�}r�>��C��!s~�~>d��χ��!���??>
���C��P�|(��>��яjй�E�s=�G=�/�{���������Çۏ��%�n�s�ׇO+�a��xK�M~񫏿ˏ��}��~��n}x�]�i���ݵ?�#�e~||���#Kp��m?���n��?|j?��x�ڭ�tw�t7������?����޼���Ǖ~\������a��o���t���P�1Y�o�ݧ���O����_{F�P>���H�����������Ut�O�s_y���7nƉ�P[=g˱e^Y��3J��£m�S�����c�[��t��xws�p��+?��|���i�}X>��� &�7%�ͻF�h�]��o�z~|?᫹p�\l�/���R�۸�G�Ekt����&]j/��6��a��=�A?;b&:Q����o�g�����KG�b}��+��x$�]��G��ǏG��ǏG��ǏG����#�������|st��u��??���[>>=����8�F������?+��O�~�p�_>�9�_%���(}e&_ĲdJ�TH-�W��必TU�zMT�`����X��*�'�9�"������8�������IP�7�L�7�˃��	�WK�U��Y��V��iU�z�����x�]���:��9s}5��@�>��+��\�"|�\$�Q��"��#�_���|D�G�Y�%I����P]>b�u&��:|jt�3	�^��e��7	g��]��c����r��؍�y�/��y�9o�O���G���t�/�r}�m�^���Ag��������g&I�k�w0]#����k8�^�k�P������}�����M�b]�ĺ��<���<����������񂮹]�6�~�>rp.�5۳�E�ey���`��������b�ݮr��I��v=��/7���_��������n��-9��-�����Ϳ��&�#M��.:=M�&A�����ᔆ���_�~���~��M����2��K��������ӏ�ڇ�W\�̳��ӷ������M�+7�N��H�ο]�?�t�S�y�!;�[s�J;��X�7G���%->��o���S�=�H���'���?O��3?������~��d��v�w�sҧ�C���5�7��%y��+Ë	l��Zp��OB>{�k�o���X����t:��������e��Ÿ�Y�p�YU�額�t���[��=���湿 �=�Ɉ���p�t��<����kI{�Z�|h1۵Ķ3����Wx�<�屓L��Z����s�}���cQ{>��]E:=6<��Wx�<����I���*}�4O"�t�&�N�濿(�%��*���t�_���_��F؛ٮ�?�.�>#���/�/O_E��vU����t1��������PK   �S����*  ��            ��    cirkitFile.jsonPK      =   +    