PK   "��S�ݚch  �_    cirkitFile.json��n�F��_����i���]�� �2�Ivn�����n�+�IAh^f�i��lK��T��c`�/�m��T�:��y��h���.��պ�خ���67�������ft�X�7��us����/�����m6]}�_-��f�T��h���N��PU6��m6We^�Ӷru;V��b�}�.m>��ec���7)
�iU�|2��s��Z�>�\=��$C�еdd+��y���YSL��q��M�ZY��m�[5�E9��J��5Y��l��9VfRL]eN��̛���|j���Z;Q�|�O�jܧW��F6w+랋
�I�����W?��l�,�W}|��k֋�?}��L
�"���K�z��{-<l����:Zx��\��	�����ӕ輩��O2z-]t�2��7��7��7��7��7��7�s�I_J�ռ�D�k�еdh��
�5��%N>�<u�C��G�V�`����cD0tߍD�A0t�i-�{�Y-�{�=q+*X7Ѳ����#����%�f�y!�!��w^H�E$C�o<���o<���P�$I~�t�8���H4��a&��q�L��zx���������`pr~�M�l�5����O�O��4�O��ܰ�V?�NSW���f�F�ks��Zӯ�ڲ�c��9�K�^.��f��w#�_��/g����,?��o_����ϱ���Һ��ѵ��ڄ���`�/X��4�O��T�����d�+Y���4�O��T�����b��X���4�O��T�����f��Y���4�O��T�t�>��!ƃ�9b)j��
�Ѹb�i���� ��6�`)0�Xu�CҰ�$��a�����U��:b���a��/��Xu��Ѱ�#��a����g��Xu��Ѱ�#��a����'(�XuإѰM#��a�����X�XuثѰY#��a���vOWvl4lو)j���)��S��U�}7b���a�*|���g`���ލ���)j��
�1�b�a���ލ���)j��
���b�������KQ�U����{7�n�5LQ�U����{7�n�5LQ�U����{7�n�5LQ���@��ލ��1ES�0E�{�R��wc`�FLQ�5LQ��K�:��ػS�0EST�W|��{7�n�5LQ_�x�j�t��j3W�y��3�M��e�l>k�.��rg�p����(�Խ������oN��LM[�����\gMn������X]ͪ�����ܓ��sO��Ͻ�n��s���ݫ�<��Veu�窘�u==�=�{?��Rsk�4�ڶ�r[�2z���R�T��\�RR���n�w�_���j-���I���/�(^��^�?��K�����E�<����k[~GIM������l�彩��_P2���[��R�� ��4Υ�1r_�Z�R"�R!(5SuP�j�)_�ԯ���S�z[�Ż��%0�*~���l�*6L��Sņ�b�T�)v��2�]���%0�*��R��߮��RE)��2Ul/Vqj:�yN�AK�853�ک�G�K/5�X݋GSj��R^��F��K�����'G���H�:Ǔ��tyW��C�������؍�<H'v� ŉ��U�81 yD����_��sspTPi�t����J����	;8*����ɣs�� ��Tg��GT�OTa���crpTP�}�<;G��H��:8*�t�͉<eG�vq'J��(=��Hy��
*��vpTP��W�����JC��HT���%yN�
*��{pTP鞯 �>8*�4D:���QI��"�?<,i�`>� �#�@�ޜU6�W6�Yƹe�e��e}_ yB<,�7�;2�ÒzCR$y��%�Ɯ�AxGR� �1�,��aI�1�lޑ�"Ho�B�~xXRo�w$∇%�ƌ� ��%�Ƽ�AxG2� �1;-��aI�1Gmޑ�$Ho�T��xXRo�W�w$g	��ւH"��s��Id��W��� ���%Y���AxG�� �1-�9�aI�1mޑ�'Ho��H�4�_�w$
��ׂ�$�����I������ d��%����AxG2� �1-�c�aI�1mޑ4*Ho�_��xXRo�_�w$�
��ׂ�'�����I������ ��%����AxG�� �1-���aI�1mޑԬ��ó ��o��Fi(��M�P.�Kj��rq]RC� �������%��a�lZi ײ}ܬ���bN䒣�^BI䒣\\��@.9
�.9���A)�
A�������^͔�f�W3��
�L	k��5SĚ�b�T����L��Sņ�b�T�a��0Ul�*�LۋU��%Ga�r�J䒣\<����(��@.9��C)9��:�x�꽼�I�`����\��hԝC���H ���� �\4*�4D:�E��J���@.T"	�QA�{.J@ �
*��rѨ��=� ��F��HG�hTP鞭�E��JC�#�\4*�t�$�E��JC�#�\4*�t�M>�E��JC�#�\4*�t�rѨ���H �
*�c��\4*�4D:�E���	f���T8,i�`>� �c�\�ޜU6�W6�Yƹe�e��e}_�\8,�7��;����fa0K�9g���r1zc�YL�Òzc�� �c�\�ޘ�Sᰤޘ�6�X �7f���T8,�7��;����ia0K�9j���r1zc�ZL�Òzc�� �c�\�ޘ�Sᰤޘ�6�X �
毅�T8,��
��;����ka0K��k���r1zs��D�@��qϤ�P�0�Z߻3D K��k���r1zc�ZL�Òzc�� �c�\�ޘ�Sᰤޘ�6�X �7毅�T8,�7��;����ka0K��k���r1zc�ZL�Òzc�� �c�\�ޘ�Sᰤޘ�6�X W��@.9��ܠ�@.9��7q���(�%9�K�rq]���(�%9�K�r8�_o�?���[�ǋ�ϣ��ތ~Z�ۇ��]3mg��r�Z������ASS)�3NL�x#��eC����l�B0�-���K�v}C'&N���i�o��{����:�Ⱥ/G2-zO4�}r>������aU�ѝd�Zt�i�F���3�L6�n�*R��@	A�����������G�o����������؍.��p' �@�! f ��g ��' �%���o�Y�O@�g�O@�u f �A<�����w�� ���g�gx[#����N菳<H�w]���|��~��|\,�c՟^��	v�돋�4q]��\Ft'�,��g���~׳oINe���t:Zr�6��Xa�<\]�E���cpE8��-crN�d�*a�ZZ{���R i�ji�n_8)@!��������Lt	�C��=yz��֩�֩�֩�֩�֩��=%'��C('x�K_X�JTua+�Qa�Ul�Tqr�z������NN_O+����jM�c�����/9�]�?r�Iܲȱ&q�"���OՑJ9đR�x��=�!�" i=�pk~�ӿ.���trt ��O�-�{�i,Y �K9�@qw�M)����!*�)F2�9<D���$�sx���nDK�'���,�؆Iz���j��%�8����"jp�r�9<DE1�Hj:����< ��b��}9	H��2���q�"��b$���CT�W ��CTS��sx���71@�9���(�	-����À�rQQL1H��1���ŏ���K �=0�X̸TK�����!,��M�д&b�A@FK1�XH8�h)�>b��  �%`��,c��R-�'��-�f���j	8=a�5�h)f�-�'��-�f��j	�<a5�h	8=0�XԶTK��	c�A@FK��Y�b��Z�O!2Z��2�-}� �}�xh�y� �}`���k����F?��������E[K�$�������|�e,�Z�%�����  �%���,c��R-�'�c-�f���j	�>a�2�h	�>0�X��TK��	c�A@FK���Y�b��Z�O�2Z��2-��}��c���}`��xg����F��������E7^�,����fI�3��%�3K����,��r������˒������[̺H��e�dҌ�~u/u�w��t����W�Î7����E��u������]���K�g귯�l�}�݇u�i�}\w��]��0]���z����z���6np�z�_�f@ڮ��r/G)/�R��å��eN��hǔ�|��;���A_S��RZ����ƾ�Ü�s�]�H��6�������H��� �l�	�a��d6������l�9���Ɉ��� ��l~���0A0i�x�� ��8S<L`��F3���w�&�����i���N_u���4�Rt3l7���q�Lڻn�pr�t��o�͛n�'-zߤ�&�o2a��7ٰ)�7�a��7����7aS�o*æj�T�M������j�p9��r�롟H됵~Z+��Isw7>�s����w��MWk��V��jn����Mָ�;i�b��B�����c3�~��f\����O>�k�n)ub���o�њ{pw�vh�F�g��0��×ͦ������֫�v�Y��ۧ�������+��Y/��<�e���k����=v?�����r�g;��z�a��_��=���{h}�C����a1�k��n��q�ng��?m���f�8o���u��?���^f�n��׏�͛�,g�]OD>+?-�Zl+��<���.�j_v�M��r��j��Ưp7�x��i}�U�֦,�:S�2����e����ui���u�,��>I7�7��'��4�����������݋�!/�[w��vo>���Vκ�<��V�F�ژݼ�s����PE��{�"��b���q�X��]?�շ�V��MZ?�UZ�jh��Mf��=:a��)���_�*�Q������f�s*+s5���c�oJW�9-�$��p֋O?l��ɬ늧��m~x���������|�T��&{�T�}M�:�m�L?{����e[y�������̙~�L?��-�MUU���m�&�]���Z��k�{��}ʪou�ܼ�}��2ǽ�ASL�}Sѷvq��M1�wMQ��M1}�M1y�M����R��o�ƾ��pR����y�We����ݶ?���x�V���ó�m+e�����͋Jeӹm���դm�f�u8�ήI�j�eٟ��ӹ��K�������G���wG ��1��9�U��lZ~|�+�Ǌ�KJ��?ְ�k(�zT==b�c���},�?������߾����w��]�y����������o�?�s�{+ݸ5�z9���:1�����\�;Ϫ��e�Z��-3��e�������^<�ۍ��>��=7�vU��w���铍��O������f�߰����O~p�R���%WJ��nċ�2�4�O������G��ں�{��ر=u�z��Yԃ=K��&�*��Nt�$:�l�s1�{���}k����߻ֵq��9�k�9q߯����l��g���/�y��K��?w*�w<l�[������k���ߦ���G���N��`P��>~���7����Y�������<����H��ܷ��ߖ��ϖ��G4ݮ���K3�w���&����W�s�?�i;��rZM]sZ�I_˞���G��,�ڽ�,k����S���,�-
�GwJ��Z����D@Z����}�6TEW�G�A}��?��PK   "��S�ݚch  �_            ��    cirkitFile.jsonPK      =   �    