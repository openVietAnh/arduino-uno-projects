PK   �S?MA�x#  S    cirkitFile.json��n�ƕ�o�P���ԩ�5���]l6	� �A���+�g[�������5m�<j5����$�x$�]�_V�K�N�p���w�n�6�������[r�Wλ��|�W{}���n��|����|����<���`�ݐ�v[�lR=6�뜱#U&dך6ԃ}CdC��&o��^������G q���}�����n�{��&�a����&t��ٛ���뜃7�\��I���J#؍i��z1k(�`7Q���B���k(�`7��A�n1�4��$1�4Bɫ��.Q(�	��!
�<I�C
i�$y�B^$��PK���dM�|I��B�s��	�S1�KYg(>io
(�b���!ay&�H�����Y�#I���_��b'Q( �ĉ:R%�H��8���*��_��J'a���)������8D��_.�!
��r!a7^n2�!
�<�C
y��(��)Q(�S�P�s�8D���Nq�B!ϝ��B�;�!
�<w�C�M��Nq�B!ϝ��B�;�!
�<w�C
��py���)Q(�S�P�s�8D���Nq�B!ϝ�v�S�P�s�8D���Nq�B!ϝ��B�;�!
�<w�C
y��(��)Q(�S�P�s�8��T��)Q(�S�P�s�,����������R
�y��ͻ�������pw�7�p��#,�-��V;(a���a�sX�t������c�����x�v����te��.b�����\��UX�t�����]��JGX:�i��>����["��#��C螰}6a�����_����G`>~��ڙ��	؛؜؝`���/��;,����T�~`���#0����T�|��w�����
���|�>0X?�c����_��vX>����`����G`>�L �9�X>��\�~`���#0Ϣ �~:�~<��?�`��ǳO�������|<o��`���3~�������|<W	��`��ǳ��������|<?��`���3��/x�����|<'��`��ǳ	�������|<��-�+Z`����Ã����|<���`��ǳf�������|<���`���3��������|<���`��ǳñ�������絃��,��xF>X?������k	���,���
X?�,�4��`����G`>�<��?�|��`����G`>����?�|��:%`����G`>����/�����|\��`���Um�������|\���`��Ǖ��������|\	�z�:z�:�D���`���#0ם��X>�q�,�~`���#0����X>�q�2�~�`������������|\��`����2%���V9�5?.ȷ��q���؈WT���l�����>W6?.Թ��q�͕͏Kc��u�^+춳�ֶv�ٲlk���l5�����y�S�шR��� ����{�����1�J�.�v���u�֯�'QoZPP��(�}�>��ׯٲNk��`���ֶ?��\����&�ܛ�z2�ȸ����K}:3�[����{J}�1B��SgRW'(��j�����/j~z�u�8�ڌ]nMp�h��l�T�Q�Cwf��{nr��X�Sg�qM]�sM����g����p�s��S�ͮqٖ�z���д��9��m
y�|���O��槏}Q�3�^c54�PHք��Mc}m�:���clCs�ؗ4?s�K��9�%�O{�c"���(8�L��hlO]{
g�}Q���N9��$2��:2M_�#��cm�rlg�������TS�+3:���ԭI�\���K����}I��{o�+]�g���K�,Y25�7>�.���������>P[W]=��B,�M6�zS�]�Œ»f8��E���:;�����\������K�/��v��g3������o��n{��]��A2^.DW����%t	hJ�(~铌�PD�(Д��~����W2"�"
(�@��	�@_~�|���(��*�F�@�o�a�@�,����Y�1�!�ӽF*���_��`y�`��N�YAL��M��[�U-d�eoe]�E��=f�)}am#�8��5���r8��8*��nk����������J�:w��,��"��:����_D�L�<��d��� &Xw�<��d� &�H����Hvz"b��q��Hvzr�aBE���,�{XGE��L0&X��<����`L�<�ay�+���`y���8*Wd�1��x��qT$�c��� ��H\�Ƅ�'��)����Q����	��,��"�,|,�XGE���(&T$��c�����H<S�����Q�xF+�	��#,��"��K,�GXGE��0&X�`y�g���`y����S��O�8���:M3CD%VRa��㉏�@]5XI��n�'D£u�`%V�9.��
�U��TX��R����FVRa-� ]�˻`�`%�2FQ����FVRa���B0�@]5XI�u6�wzk����q�xT��������ǥBK:��n���J�K�v��.�1^��ThI���5��V�}�В-�3����S�%Z~�_G[�BK:�<�AG['�BK:�<CG[7�BK:�<�DG[G�BK:�<7FG[W�BK:�<�G����/S�%Z������/S�%Z�s����1�Gb:����2���ThI�����h���ThI�����h���ThI���$�h���ThI���V�h���ThI����h���ThI����h���ThI����꼘���ThI����h���ThI���P�h���ThI����h������:����2���ThI�����h���ThI��k�h���ThI��k%�h���ThI��k>�h���ThI��kW�h���ThI��kp�ht|�
-��r-mu|�
-��rMmu|�
-��rmmu|�
-��r�m�f�)M%��eAǗ_�BK:�\3HG[_�BK:�\�HG[_�BK:�\�IG[_�BK:�\�JG[_�BK:�\SKEۨ��ThI��k��h���ThI��k��h���ThI��k��h���ThI��k��h���ThI��k��h�T�C�̇�/�:�,��2Zҡ�Z�:���2Zҡ嚌:���2Zҡ�ڒ:���2Zҡ��*�V:�L��th�֧��:�L��th�f���:�L����>�������.�����1{3t>u}�sp�u�WF9Q�ve��dWF9Q�{e�k\��r�V��('�[��r���('*H��r����^꼘�{j�׵a0���Ҫk�`z�P׆�����0O��x���a�^<_V}mֳ��:^y|mP���S�T�3���·k��{�lֵa���:^tmL&>�H��0�\|j)µa.�����}o�ͽ	�'���������ԧˣ�EQ.����hc06�rH}�L��d�PUm���̲(�E��m��]m�.�&�\��m6}*�����,��\d�M��`�cK�L3���kr�)�����,��`X.&�EQ.�<�]�-��2�7�ik�r&�m
y���ˢ(uY�.��\֥�jh����	cߛ���tutm��؆f�.K�\�eI�˺,�rQ�6�D.:��mp֙����>��6�.�(�E](甚D�*�Ȅ֑i��֘�kە�̲(�e�j�reFG����5)�<�XG_�ż�eI��,mt���l\}��%q������å��~��^�"�@m]u�X.cE��7��n�M�w}�5�k��,��\λv,=�&��d[�ٗ/D�|���.vy�5`I�C��0�����!?Wox�~��v���o�J9�@��!�_# D�@����Nw� D�@v�3!��].(���A�@��t�B
d�;y"P ��+�I����K۰�M�č�d�7?1L��M�䍊d��e1L��M���d�7�1L�N�$��d���1L�<�`y��o�c�p�o� ��,��"���,�;XGE���&Xw�<��d��_0L�<�`y��a�8,�{XGE�j0&ܝܭX��<��ĵ�`L�<�ay�k-��`y���8*���1��x��qT$�%c��� ��H\�Ƅ�'��)����Q����	��,��"qM,�XGE�9��G?�<ay��lØ`y<��8*��1�n�o��x��qT$��	c�����H<w���,��"�\5,�W�<~*��yg�y����a����J*�v3�ӈ�
�U��TX�f6���+���ͬ�:*PWVRa-�KE�Yy����Z�A*��J�@�`%�2FQ�uVV��+���ͬ�:*PWVRa��Y=tT�����j7�Z2�@]5XI���	�1:�K��th��fm�\�����]�c�H�y�В-�k�����R�%Z~g^G[�BK:���:.L��thy���:NL��thy.���:nL��thyN���:�L��thyn���:�L��thy��΃_�BK:�<WIG[_�BK:�<�JG[�'bJ��t|���eNǗ�В-ρ��VǗ�В-����VǗ�В-�I��VǗ�В-ϭ��VǗ�В-���VǗ�В-�u��VǗ�В-���y1IǗ�В-�=��VǗ�В-ϡ��VǗ�В-���V�mE��u|���e^Ǘ�В-����VǗ�В-���VǗ�В-�J��VǗ�В-�|��VǗ�В-׮��VǗ�В-��P�6��2Zҡ�Z":���2Zҡ�(:���2Zҡ��.:���2Zҡ�5:�*�$S�J��˂�/:�L��th�f���:�L��th�����:�L��th�����:�L��th����:�L��th�����QǗ�В-���VǗ�В-�8��VǗ�В-�j��VǗ�В-ל��VǗ�В-����V�ʇR�_u|Y��e*��C˵u���e*��C�5u���e*��C˵%u���e*��C�52U��t|�
-��r�Omu|�
-��r�Rmu|�
--�}^*:6)��Me]0���ic�f�|��:���S�0��r�6��('�ɮ�r����('*o��r�V��('�[��r���('*H��r����^꼘�{j�׵a0���Ҫk�`z�L׆���S˄���ŧ�\��1���*�k�`z� ׆���S+.���ŧ�5\{����S�>��\����&�ܛ�z2�ȸ����K}�<�Y�"KO��6cC(�ԧΤ�N&PU�V���,��\d���y��f�rk��E��fӧrL��͡�̲(�E���86�1��D��4�8��&�2�͝�̲(
��b�[�bγ�5.�2�/�z��6y g���M!c��uY�.��\�eQ�˺T�XM4�5a�{�X_����m���,�eI�˺,�rY�%Q.����Eg����:Ӷ6���S�ƞ�e]E���R��Td���L������Xۮ�e�EQ.��TS�+3:���խI�����:���(�,K�\di�+��g���K�.�;5�7>�.���\��(Yj몫�r+����&wCo��X�1]3\fY�r޵c�im0��%3��5Ⱦ|!B���v��K�K���x]����M����67�_����W������[>����f����ۯ�~��G�-mE��]���}�RB�AF Ԁ3ʼ�t�I�I��/VM�e��_���{�2�.�{���{_Dt���Q�w?e��������]�Z���@���O���z9T����"qq� ��
�B!�bb����	��^?!���+�)_O��7w���C~�7����8���y�no���?H�c�d����h�/�2(�C9�4���^G�D��C�4�vz0~$M%��r�J.�8����)�!���_H!a����v���C��_T�r �+ҫ<�ݿ*!� ���]��l&�!�)��Dİ��?��\bb���H�ȼ�v�v��#�%v2��m�Ys��� �Y��_ߑr���^����v�>���� 5�c��MR�����v�N���| ��c��[]By�-L�H��^�1�F0��O= ��cp�Y  �z@>����� @>��|*���2�| �T�k08 �4 �<��p n�"���i �Sy��� �� ȧ�\��ȧ�O�1���C�k'8 �4�<��p �i�Sy��� ��ȧ�\C�ȧ�O�1�6��O+@>���� @>� �tc�k&�:�x�B�x�#0���j]��A�����nf�,p� �a��g7�Z��x��|�+~�߬P��x�|�+��~�b�����������
�	��G`>�����Ń��#0��5���y�[�9g��x9g%�p� �a���/D���hC&$4!�̉�nJ�mK�KmL���&�h���	��Є�0ZC�A���VFk�6)`BB��h�FLHhB~-�!ڬ�		M�ﰣ5D;0!�	��{��h�&$4!O@߷F�0!�	yfZC�O��ge�5�?@�?AA���)�S���&��/h�>LHhB�����S���&�iGh�>LHhB�2���S���&��^h�>LHhB�����S���&�iv��C�>LHhB�"���S���&��h�>LHhB�������m/�O�h���>LHhB����S���&��h�>LHhB�����S���&�i�h�>LHhB����S���&���`ڧ�		M�S���}
��Є\6 �!ڧ�		M�%��}
��Є\��!|b
|f
ڧ�O	h�&$4!��@k��)`BBr���h�&$4!�'Ak��)`BBri��h�&$4!��k�>LHhB.i���S���&�r<h�>LHhB.%���S���&�2Hh�>LHhB.��>�>��S"ڧD�O��Kg�5D�0!�	��ZC�O��K��5D�0!�	��X�
�S���&�Rqh�>LHhB.s���S��t�p�2����k�����\�~Vju����YnV�te�Y�ҕ�g�EW��U]�~V�smw�Gi��/�6��K�WP[@��랭_��|�����_�u�:��8]����UA���Ui/��Y�~���ޭ_J���l��>�V��x��;_}im i�w�6��n[�޵��M��7!�dR5�quUu!x��tn4��������hc06�r }�L��d�PUm��?��E���n�}W��˭	.s�M���6�����?����86�1�����4�8��&�2�̝?��E��?���?��lv�˶���Xڄ��MșP��m
y�+��l���?s��ڟ;�j����B�&�}o�k��ѵmc��ǿ����_����/i�����L7�V�Yg��Fc�8x���S8w��ڟ9~�9�&����֑i��Ę�kە�;��E���ߦ��\��Q,��nM��]6�ї�D1�����g��FWz����ї�YRgj\o|.?\[�Ϻ�E�������z,��Z�lr7���%�w�pn��ڟ�v,}�&��|m��ٗ�*_Ҹ�b����%��������M�y�nJ����?\-��_����=0��x�ţ"l� ��<�o��f� ���ğ%�0�?N�y��-�pSlnḅ��[8nḅ��[xnQ������K�%W��\f_4Xr]�+Z.I�7\�	_m�$��8�%9�e�I�E�%���|_��ߛ��������ٔ�,��=���÷���𾖴w��TA���I悐H�i�t�ל9)Q���9�9�ߝi7��әE!����>��@»Js�����r��#G�v�����mn�[N��ly����3NZ�1m��&����7��M~�)<m
�M�iS�o��6U�M�Ӧ��U��vs�	n��������O�"�br7�=�����tć��3��5?�E���O��m����a~���po(Gy������(p����y���w����դ�xwS�ʿ�����ww���Wo�|{?�����O7�7����o��ov<�z(�E�o��㘻��ݰ;p���]�xs���ҏon�E������:v����ob��	��4+־��zS�ц���L.�Ӵ����u�a�x�!�u�6�F��W��M9_yOs�������u���,��{�Sc�]3m}�K<�����-�`��-Tn	���Ï��{��9�P�����R�8����{�ť�-e�}�Ku�%n�[�p�=ز?��~���/�p�?�B�[����`C����M��n�zx�o�v���Ho�*�C�������+�����n��r8�/` ������@�W<׋�^q��b����@���jF3�vh��*7��߽E�q�w/L=�d>����������ޓ'�ˣs>V�XW��ˤ좩�(�u����/��KN�oN����'?N�O��O~<>�!=�W����O�7��g�z?��IC����4��q/XtOgQ/��
؛t�_�:Ex��lV�#���WU�_���H�g����������g���;^\m?��T_�r��y�ӋkG�Jwi�/#�J�2)=���ڔ�㎳��ޒ����^�����q�i��h��fO���>�5��V�����(�b��/�b��u�W��ȶ\�޼4������>u2�Nf�ڢGKz[s215����S��	���0�����4��G>N���>�dg�����stf���ĩ�M��|�?v���ښRr1���D|����awLS����w�<ϟz�s�|6�󉸟R�qӟʡ�L�M�v��_�/��+�r��������w�g��w��Y���P����/�����>�"�\G��q��kW�j,&��ٗQ}��e��!�]��|��=�:���m��r{�
/}䭀O=��c�}r��N��Q�N��z�O����Ϫ_F7��@�t�����4v�Wx?�؟S�ݻ`��~�+%�:�Ӄw���S��y�˽s�~y0�#i]���>�jE�S����¾ӧ�����х5ar좗����`����
�������PK   �S?MA�x#  S            ��    cirkitFile.jsonPK      =   �#    